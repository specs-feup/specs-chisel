module SCIEPipelined #(parameter XLEN = 32)(
  input         clock,
  input         reset,
  input         valid,
  input  [31:0] insn,
  input  [31:0] rs1,
  input  [31:0] rs2,
  output [31:0] rd
);
  reg [31:0] coeffs_0;
  reg [31:0] coeffs_1;
  reg [31:0] coeffs_2;
  reg [31:0] coeffs_3;
  reg [31:0] coeffs_4;
  reg [31:0] coeffs_5;
  reg [31:0] coeffs_6;
  reg [31:0] coeffs_7;
  reg [31:0] coeffs_8;
  reg [31:0] coeffs_9;
  reg [31:0] coeffs_10;
  reg [31:0] coeffs_11;
  reg [31:0] coeffs_12;
  reg [31:0] coeffs_13;
  reg [31:0] coeffs_14;
  reg [31:0] coeffs_15;
  reg [31:0] coeffs_16;
  reg [31:0] coeffs_17;
  reg [31:0] coeffs_18;
  reg [31:0] coeffs_19;
  reg [31:0] coeffs_20;
  reg [31:0] coeffs_21;
  reg [31:0] coeffs_22;
  reg [31:0] coeffs_23;
  reg [31:0] coeffs_24;
  reg [31:0] coeffs_25;
  reg [31:0] coeffs_26;
  reg [31:0] coeffs_27;
  reg [31:0] coeffs_28;
  reg [31:0] coeffs_29;
  reg [31:0] coeffs_30;
  reg [31:0] coeffs_31;
  reg [31:0] coeffs_32;
  reg [31:0] coeffs_33;
  reg [31:0] coeffs_34;
  reg [31:0] coeffs_35;
  reg [31:0] coeffs_36;
  reg [31:0] coeffs_37;
  reg [31:0] coeffs_38;
  reg [31:0] coeffs_39;
  reg [31:0] coeffs_40;
  reg [31:0] coeffs_41;
  reg [31:0] coeffs_42;
  reg [31:0] coeffs_43;
  reg [31:0] coeffs_44;
  reg [31:0] coeffs_45;
  reg [31:0] coeffs_46;
  reg [31:0] coeffs_47;
  reg [31:0] coeffs_48;
  reg [31:0] coeffs_49;
  reg [31:0] coeffs_50;
  reg [31:0] coeffs_51;
  reg [31:0] coeffs_52;
  reg [31:0] coeffs_53;
  reg [31:0] coeffs_54;
  reg [31:0] coeffs_55;
  reg [31:0] coeffs_56;
  reg [31:0] coeffs_57;
  reg [31:0] coeffs_58;
  reg [31:0] coeffs_59;
  reg [31:0] coeffs_60;
  reg [31:0] coeffs_61;
  reg [31:0] coeffs_62;
  reg [31:0] coeffs_63;
  reg [31:0] coeffs_64;
  reg [31:0] coeffs_65;
  reg [31:0] coeffs_66;
  reg [31:0] coeffs_67;
  reg [31:0] coeffs_68;
  reg [31:0] coeffs_69;
  reg [31:0] coeffs_70;
  reg [31:0] coeffs_71;
  reg [31:0] coeffs_72;
  reg [31:0] coeffs_73;
  reg [31:0] coeffs_74;
  reg [31:0] coeffs_75;
  reg [31:0] coeffs_76;
  reg [31:0] coeffs_77;
  reg [31:0] coeffs_78;
  reg [31:0] coeffs_79;
  reg [31:0] coeffs_80;
  reg [31:0] coeffs_81;
  reg [31:0] coeffs_82;
  reg [31:0] coeffs_83;
  reg [31:0] coeffs_84;
  reg [31:0] coeffs_85;
  reg [31:0] coeffs_86;
  reg [31:0] coeffs_87;
  reg [31:0] coeffs_88;
  reg [31:0] coeffs_89;
  reg [31:0] coeffs_90;
  reg [31:0] coeffs_91;
  reg [31:0] coeffs_92;
  reg [31:0] coeffs_93;
  reg [31:0] coeffs_94;
  reg [31:0] coeffs_95;
  reg [31:0] coeffs_96;
  reg [31:0] coeffs_97;
  reg [31:0] coeffs_98;
  reg [31:0] coeffs_99;
  reg [31:0] coeffs_100;
  reg [31:0] coeffs_101;
  reg [31:0] coeffs_102;
  reg [31:0] coeffs_103;
  reg [31:0] coeffs_104;
  reg [31:0] coeffs_105;
  reg [31:0] coeffs_106;
  reg [31:0] coeffs_107;
  reg [31:0] coeffs_108;
  reg [31:0] coeffs_109;
  reg [31:0] coeffs_110;
  reg [31:0] coeffs_111;
  reg [31:0] coeffs_112;
  reg [31:0] coeffs_113;
  reg [31:0] coeffs_114;
  reg [31:0] coeffs_115;
  reg [31:0] coeffs_116;
  reg [31:0] coeffs_117;
  reg [31:0] coeffs_118;
  reg [31:0] coeffs_119;
  reg [31:0] coeffs_120;
  reg [31:0] coeffs_121;
  reg [31:0] coeffs_122;
  reg [31:0] coeffs_123;
  reg [31:0] coeffs_124;
  reg [31:0] coeffs_125;
  reg [31:0] coeffs_126;
  reg [31:0] coeffs_127;
  reg [31:0] coeffs_128;
  reg [31:0] coeffs_129;
  reg [31:0] coeffs_130;
  reg [31:0] coeffs_131;
  reg [31:0] coeffs_132;
  reg [31:0] coeffs_133;
  reg [31:0] coeffs_134;
  reg [31:0] coeffs_135;
  reg [31:0] coeffs_136;
  reg [31:0] coeffs_137;
  reg [31:0] coeffs_138;
  reg [31:0] coeffs_139;
  reg [31:0] coeffs_140;
  reg [31:0] coeffs_141;
  reg [31:0] coeffs_142;
  reg [31:0] coeffs_143;
  reg [31:0] coeffs_144;
  reg [31:0] coeffs_145;
  reg [31:0] coeffs_146;
  reg [31:0] coeffs_147;
  reg [31:0] coeffs_148;
  reg [31:0] coeffs_149;
  reg [31:0] coeffs_150;
  reg [31:0] coeffs_151;
  reg [31:0] coeffs_152;
  reg [31:0] coeffs_153;
  reg [31:0] coeffs_154;
  reg [31:0] coeffs_155;
  reg [31:0] coeffs_156;
  reg [31:0] coeffs_157;
  reg [31:0] coeffs_158;
  reg [31:0] coeffs_159;
  reg [31:0] coeffs_160;
  reg [31:0] coeffs_161;
  reg [31:0] coeffs_162;
  reg [31:0] coeffs_163;
  reg [31:0] coeffs_164;
  reg [31:0] coeffs_165;
  reg [31:0] coeffs_166;
  reg [31:0] coeffs_167;
  reg [31:0] coeffs_168;
  reg [31:0] coeffs_169;
  reg [31:0] coeffs_170;
  reg [31:0] coeffs_171;
  reg [31:0] coeffs_172;
  reg [31:0] coeffs_173;
  reg [31:0] coeffs_174;
  reg [31:0] coeffs_175;
  reg [31:0] coeffs_176;
  reg [31:0] coeffs_177;
  reg [31:0] coeffs_178;
  reg [31:0] coeffs_179;
  reg [31:0] coeffs_180;
  reg [31:0] coeffs_181;
  reg [31:0] coeffs_182;
  reg [31:0] coeffs_183;
  reg [31:0] coeffs_184;
  reg [31:0] coeffs_185;
  reg [31:0] coeffs_186;
  reg [31:0] coeffs_187;
  reg [31:0] coeffs_188;
  reg [31:0] coeffs_189;
  reg [31:0] coeffs_190;
  reg [31:0] coeffs_191;
  reg [31:0] coeffs_192;
  reg [31:0] coeffs_193;
  reg [31:0] coeffs_194;
  reg [31:0] coeffs_195;
  reg [31:0] coeffs_196;
  reg [31:0] coeffs_197;
  reg [31:0] coeffs_198;
  reg [31:0] coeffs_199;
  reg [31:0] data_0;
  reg [31:0] data_1;
  reg [31:0] data_2;
  reg [31:0] data_3;
  reg [31:0] data_4;
  reg [31:0] data_5;
  reg [31:0] data_6;
  reg [31:0] data_7;
  reg [31:0] data_8;
  reg [31:0] data_9;
  reg [31:0] data_10;
  reg [31:0] data_11;
  reg [31:0] data_12;
  reg [31:0] data_13;
  reg [31:0] data_14;
  reg [31:0] data_15;
  reg [31:0] data_16;
  reg [31:0] data_17;
  reg [31:0] data_18;
  reg [31:0] data_19;
  reg [31:0] data_20;
  reg [31:0] data_21;
  reg [31:0] data_22;
  reg [31:0] data_23;
  reg [31:0] data_24;
  reg [31:0] data_25;
  reg [31:0] data_26;
  reg [31:0] data_27;
  reg [31:0] data_28;
  reg [31:0] data_29;
  reg [31:0] data_30;
  reg [31:0] data_31;
  reg [31:0] data_32;
  reg [31:0] data_33;
  reg [31:0] data_34;
  reg [31:0] data_35;
  reg [31:0] data_36;
  reg [31:0] data_37;
  reg [31:0] data_38;
  reg [31:0] data_39;
  reg [31:0] data_40;
  reg [31:0] data_41;
  reg [31:0] data_42;
  reg [31:0] data_43;
  reg [31:0] data_44;
  reg [31:0] data_45;
  reg [31:0] data_46;
  reg [31:0] data_47;
  reg [31:0] data_48;
  reg [31:0] data_49;
  reg [31:0] data_50;
  reg [31:0] data_51;
  reg [31:0] data_52;
  reg [31:0] data_53;
  reg [31:0] data_54;
  reg [31:0] data_55;
  reg [31:0] data_56;
  reg [31:0] data_57;
  reg [31:0] data_58;
  reg [31:0] data_59;
  reg [31:0] data_60;
  reg [31:0] data_61;
  reg [31:0] data_62;
  reg [31:0] data_63;
  reg [31:0] data_64;
  reg [31:0] data_65;
  reg [31:0] data_66;
  reg [31:0] data_67;
  reg [31:0] data_68;
  reg [31:0] data_69;
  reg [31:0] data_70;
  reg [31:0] data_71;
  reg [31:0] data_72;
  reg [31:0] data_73;
  reg [31:0] data_74;
  reg [31:0] data_75;
  reg [31:0] data_76;
  reg [31:0] data_77;
  reg [31:0] data_78;
  reg [31:0] data_79;
  reg [31:0] data_80;
  reg [31:0] data_81;
  reg [31:0] data_82;
  reg [31:0] data_83;
  reg [31:0] data_84;
  reg [31:0] data_85;
  reg [31:0] data_86;
  reg [31:0] data_87;
  reg [31:0] data_88;
  reg [31:0] data_89;
  reg [31:0] data_90;
  reg [31:0] data_91;
  reg [31:0] data_92;
  reg [31:0] data_93;
  reg [31:0] data_94;
  reg [31:0] data_95;
  reg [31:0] data_96;
  reg [31:0] data_97;
  reg [31:0] data_98;
  reg [31:0] data_99;
  reg [31:0] data_100;
  reg [31:0] data_101;
  reg [31:0] data_102;
  reg [31:0] data_103;
  reg [31:0] data_104;
  reg [31:0] data_105;
  reg [31:0] data_106;
  reg [31:0] data_107;
  reg [31:0] data_108;
  reg [31:0] data_109;
  reg [31:0] data_110;
  reg [31:0] data_111;
  reg [31:0] data_112;
  reg [31:0] data_113;
  reg [31:0] data_114;
  reg [31:0] data_115;
  reg [31:0] data_116;
  reg [31:0] data_117;
  reg [31:0] data_118;
  reg [31:0] data_119;
  reg [31:0] data_120;
  reg [31:0] data_121;
  reg [31:0] data_122;
  reg [31:0] data_123;
  reg [31:0] data_124;
  reg [31:0] data_125;
  reg [31:0] data_126;
  reg [31:0] data_127;
  reg [31:0] data_128;
  reg [31:0] data_129;
  reg [31:0] data_130;
  reg [31:0] data_131;
  reg [31:0] data_132;
  reg [31:0] data_133;
  reg [31:0] data_134;
  reg [31:0] data_135;
  reg [31:0] data_136;
  reg [31:0] data_137;
  reg [31:0] data_138;
  reg [31:0] data_139;
  reg [31:0] data_140;
  reg [31:0] data_141;
  reg [31:0] data_142;
  reg [31:0] data_143;
  reg [31:0] data_144;
  reg [31:0] data_145;
  reg [31:0] data_146;
  reg [31:0] data_147;
  reg [31:0] data_148;
  reg [31:0] data_149;
  reg [31:0] data_150;
  reg [31:0] data_151;
  reg [31:0] data_152;
  reg [31:0] data_153;
  reg [31:0] data_154;
  reg [31:0] data_155;
  reg [31:0] data_156;
  reg [31:0] data_157;
  reg [31:0] data_158;
  reg [31:0] data_159;
  reg [31:0] data_160;
  reg [31:0] data_161;
  reg [31:0] data_162;
  reg [31:0] data_163;
  reg [31:0] data_164;
  reg [31:0] data_165;
  reg [31:0] data_166;
  reg [31:0] data_167;
  reg [31:0] data_168;
  reg [31:0] data_169;
  reg [31:0] data_170;
  reg [31:0] data_171;
  reg [31:0] data_172;
  reg [31:0] data_173;
  reg [31:0] data_174;
  reg [31:0] data_175;
  reg [31:0] data_176;
  reg [31:0] data_177;
  reg [31:0] data_178;
  reg [31:0] data_179;
  reg [31:0] data_180;
  reg [31:0] data_181;
  reg [31:0] data_182;
  reg [31:0] data_183;
  reg [31:0] data_184;
  reg [31:0] data_185;
  reg [31:0] data_186;
  reg [31:0] data_187;
  reg [31:0] data_188;
  reg [31:0] data_189;
  reg [31:0] data_190;
  reg [31:0] data_191;
  reg [31:0] data_192;
  reg [31:0] data_193;
  reg [31:0] data_194;
  reg [31:0] data_195;
  reg [31:0] data_196;
  reg [31:0] data_197;
  reg [31:0] data_198;
  reg [31:0] data_199;
  reg [63:0] result;
  wire [31:0] _GEN_201 = 8'h1 == rs2[7:0] ? $signed(coeffs_1) : $signed(coeffs_0);
  wire [31:0] _GEN_202 = 8'h2 == rs2[7:0] ? $signed(coeffs_2) : $signed(_GEN_201);
  wire [31:0] _GEN_203 = 8'h3 == rs2[7:0] ? $signed(coeffs_3) : $signed(_GEN_202);
  wire [31:0] _GEN_204 = 8'h4 == rs2[7:0] ? $signed(coeffs_4) : $signed(_GEN_203);
  wire [31:0] _GEN_205 = 8'h5 == rs2[7:0] ? $signed(coeffs_5) : $signed(_GEN_204);
  wire [31:0] _GEN_206 = 8'h6 == rs2[7:0] ? $signed(coeffs_6) : $signed(_GEN_205);
  wire [31:0] _GEN_207 = 8'h7 == rs2[7:0] ? $signed(coeffs_7) : $signed(_GEN_206);
  wire [31:0] _GEN_208 = 8'h8 == rs2[7:0] ? $signed(coeffs_8) : $signed(_GEN_207);
  wire [31:0] _GEN_209 = 8'h9 == rs2[7:0] ? $signed(coeffs_9) : $signed(_GEN_208);
  wire [31:0] _GEN_210 = 8'ha == rs2[7:0] ? $signed(coeffs_10) : $signed(_GEN_209);
  wire [31:0] _GEN_211 = 8'hb == rs2[7:0] ? $signed(coeffs_11) : $signed(_GEN_210);
  wire [31:0] _GEN_212 = 8'hc == rs2[7:0] ? $signed(coeffs_12) : $signed(_GEN_211);
  wire [31:0] _GEN_213 = 8'hd == rs2[7:0] ? $signed(coeffs_13) : $signed(_GEN_212);
  wire [31:0] _GEN_214 = 8'he == rs2[7:0] ? $signed(coeffs_14) : $signed(_GEN_213);
  wire [31:0] _GEN_215 = 8'hf == rs2[7:0] ? $signed(coeffs_15) : $signed(_GEN_214);
  wire [31:0] _GEN_216 = 8'h10 == rs2[7:0] ? $signed(coeffs_16) : $signed(_GEN_215);
  wire [31:0] _GEN_217 = 8'h11 == rs2[7:0] ? $signed(coeffs_17) : $signed(_GEN_216);
  wire [31:0] _GEN_218 = 8'h12 == rs2[7:0] ? $signed(coeffs_18) : $signed(_GEN_217);
  wire [31:0] _GEN_219 = 8'h13 == rs2[7:0] ? $signed(coeffs_19) : $signed(_GEN_218);
  wire [31:0] _GEN_220 = 8'h14 == rs2[7:0] ? $signed(coeffs_20) : $signed(_GEN_219);
  wire [31:0] _GEN_221 = 8'h15 == rs2[7:0] ? $signed(coeffs_21) : $signed(_GEN_220);
  wire [31:0] _GEN_222 = 8'h16 == rs2[7:0] ? $signed(coeffs_22) : $signed(_GEN_221);
  wire [31:0] _GEN_223 = 8'h17 == rs2[7:0] ? $signed(coeffs_23) : $signed(_GEN_222);
  wire [31:0] _GEN_224 = 8'h18 == rs2[7:0] ? $signed(coeffs_24) : $signed(_GEN_223);
  wire [31:0] _GEN_225 = 8'h19 == rs2[7:0] ? $signed(coeffs_25) : $signed(_GEN_224);
  wire [31:0] _GEN_226 = 8'h1a == rs2[7:0] ? $signed(coeffs_26) : $signed(_GEN_225);
  wire [31:0] _GEN_227 = 8'h1b == rs2[7:0] ? $signed(coeffs_27) : $signed(_GEN_226);
  wire [31:0] _GEN_228 = 8'h1c == rs2[7:0] ? $signed(coeffs_28) : $signed(_GEN_227);
  wire [31:0] _GEN_229 = 8'h1d == rs2[7:0] ? $signed(coeffs_29) : $signed(_GEN_228);
  wire [31:0] _GEN_230 = 8'h1e == rs2[7:0] ? $signed(coeffs_30) : $signed(_GEN_229);
  wire [31:0] _GEN_231 = 8'h1f == rs2[7:0] ? $signed(coeffs_31) : $signed(_GEN_230);
  wire [31:0] _GEN_232 = 8'h20 == rs2[7:0] ? $signed(coeffs_32) : $signed(_GEN_231);
  wire [31:0] _GEN_233 = 8'h21 == rs2[7:0] ? $signed(coeffs_33) : $signed(_GEN_232);
  wire [31:0] _GEN_234 = 8'h22 == rs2[7:0] ? $signed(coeffs_34) : $signed(_GEN_233);
  wire [31:0] _GEN_235 = 8'h23 == rs2[7:0] ? $signed(coeffs_35) : $signed(_GEN_234);
  wire [31:0] _GEN_236 = 8'h24 == rs2[7:0] ? $signed(coeffs_36) : $signed(_GEN_235);
  wire [31:0] _GEN_237 = 8'h25 == rs2[7:0] ? $signed(coeffs_37) : $signed(_GEN_236);
  wire [31:0] _GEN_238 = 8'h26 == rs2[7:0] ? $signed(coeffs_38) : $signed(_GEN_237);
  wire [31:0] _GEN_239 = 8'h27 == rs2[7:0] ? $signed(coeffs_39) : $signed(_GEN_238);
  wire [31:0] _GEN_240 = 8'h28 == rs2[7:0] ? $signed(coeffs_40) : $signed(_GEN_239);
  wire [31:0] _GEN_241 = 8'h29 == rs2[7:0] ? $signed(coeffs_41) : $signed(_GEN_240);
  wire [31:0] _GEN_242 = 8'h2a == rs2[7:0] ? $signed(coeffs_42) : $signed(_GEN_241);
  wire [31:0] _GEN_243 = 8'h2b == rs2[7:0] ? $signed(coeffs_43) : $signed(_GEN_242);
  wire [31:0] _GEN_244 = 8'h2c == rs2[7:0] ? $signed(coeffs_44) : $signed(_GEN_243);
  wire [31:0] _GEN_245 = 8'h2d == rs2[7:0] ? $signed(coeffs_45) : $signed(_GEN_244);
  wire [31:0] _GEN_246 = 8'h2e == rs2[7:0] ? $signed(coeffs_46) : $signed(_GEN_245);
  wire [31:0] _GEN_247 = 8'h2f == rs2[7:0] ? $signed(coeffs_47) : $signed(_GEN_246);
  wire [31:0] _GEN_248 = 8'h30 == rs2[7:0] ? $signed(coeffs_48) : $signed(_GEN_247);
  wire [31:0] _GEN_249 = 8'h31 == rs2[7:0] ? $signed(coeffs_49) : $signed(_GEN_248);
  wire [31:0] _GEN_250 = 8'h32 == rs2[7:0] ? $signed(coeffs_50) : $signed(_GEN_249);
  wire [31:0] _GEN_251 = 8'h33 == rs2[7:0] ? $signed(coeffs_51) : $signed(_GEN_250);
  wire [31:0] _GEN_252 = 8'h34 == rs2[7:0] ? $signed(coeffs_52) : $signed(_GEN_251);
  wire [31:0] _GEN_253 = 8'h35 == rs2[7:0] ? $signed(coeffs_53) : $signed(_GEN_252);
  wire [31:0] _GEN_254 = 8'h36 == rs2[7:0] ? $signed(coeffs_54) : $signed(_GEN_253);
  wire [31:0] _GEN_255 = 8'h37 == rs2[7:0] ? $signed(coeffs_55) : $signed(_GEN_254);
  wire [31:0] _GEN_256 = 8'h38 == rs2[7:0] ? $signed(coeffs_56) : $signed(_GEN_255);
  wire [31:0] _GEN_257 = 8'h39 == rs2[7:0] ? $signed(coeffs_57) : $signed(_GEN_256);
  wire [31:0] _GEN_258 = 8'h3a == rs2[7:0] ? $signed(coeffs_58) : $signed(_GEN_257);
  wire [31:0] _GEN_259 = 8'h3b == rs2[7:0] ? $signed(coeffs_59) : $signed(_GEN_258);
  wire [31:0] _GEN_260 = 8'h3c == rs2[7:0] ? $signed(coeffs_60) : $signed(_GEN_259);
  wire [31:0] _GEN_261 = 8'h3d == rs2[7:0] ? $signed(coeffs_61) : $signed(_GEN_260);
  wire [31:0] _GEN_262 = 8'h3e == rs2[7:0] ? $signed(coeffs_62) : $signed(_GEN_261);
  wire [31:0] _GEN_263 = 8'h3f == rs2[7:0] ? $signed(coeffs_63) : $signed(_GEN_262);
  wire [31:0] _GEN_264 = 8'h40 == rs2[7:0] ? $signed(coeffs_64) : $signed(_GEN_263);
  wire [31:0] _GEN_265 = 8'h41 == rs2[7:0] ? $signed(coeffs_65) : $signed(_GEN_264);
  wire [31:0] _GEN_266 = 8'h42 == rs2[7:0] ? $signed(coeffs_66) : $signed(_GEN_265);
  wire [31:0] _GEN_267 = 8'h43 == rs2[7:0] ? $signed(coeffs_67) : $signed(_GEN_266);
  wire [31:0] _GEN_268 = 8'h44 == rs2[7:0] ? $signed(coeffs_68) : $signed(_GEN_267);
  wire [31:0] _GEN_269 = 8'h45 == rs2[7:0] ? $signed(coeffs_69) : $signed(_GEN_268);
  wire [31:0] _GEN_270 = 8'h46 == rs2[7:0] ? $signed(coeffs_70) : $signed(_GEN_269);
  wire [31:0] _GEN_271 = 8'h47 == rs2[7:0] ? $signed(coeffs_71) : $signed(_GEN_270);
  wire [31:0] _GEN_272 = 8'h48 == rs2[7:0] ? $signed(coeffs_72) : $signed(_GEN_271);
  wire [31:0] _GEN_273 = 8'h49 == rs2[7:0] ? $signed(coeffs_73) : $signed(_GEN_272);
  wire [31:0] _GEN_274 = 8'h4a == rs2[7:0] ? $signed(coeffs_74) : $signed(_GEN_273);
  wire [31:0] _GEN_275 = 8'h4b == rs2[7:0] ? $signed(coeffs_75) : $signed(_GEN_274);
  wire [31:0] _GEN_276 = 8'h4c == rs2[7:0] ? $signed(coeffs_76) : $signed(_GEN_275);
  wire [31:0] _GEN_277 = 8'h4d == rs2[7:0] ? $signed(coeffs_77) : $signed(_GEN_276);
  wire [31:0] _GEN_278 = 8'h4e == rs2[7:0] ? $signed(coeffs_78) : $signed(_GEN_277);
  wire [31:0] _GEN_279 = 8'h4f == rs2[7:0] ? $signed(coeffs_79) : $signed(_GEN_278);
  wire [31:0] _GEN_280 = 8'h50 == rs2[7:0] ? $signed(coeffs_80) : $signed(_GEN_279);
  wire [31:0] _GEN_281 = 8'h51 == rs2[7:0] ? $signed(coeffs_81) : $signed(_GEN_280);
  wire [31:0] _GEN_282 = 8'h52 == rs2[7:0] ? $signed(coeffs_82) : $signed(_GEN_281);
  wire [31:0] _GEN_283 = 8'h53 == rs2[7:0] ? $signed(coeffs_83) : $signed(_GEN_282);
  wire [31:0] _GEN_284 = 8'h54 == rs2[7:0] ? $signed(coeffs_84) : $signed(_GEN_283);
  wire [31:0] _GEN_285 = 8'h55 == rs2[7:0] ? $signed(coeffs_85) : $signed(_GEN_284);
  wire [31:0] _GEN_286 = 8'h56 == rs2[7:0] ? $signed(coeffs_86) : $signed(_GEN_285);
  wire [31:0] _GEN_287 = 8'h57 == rs2[7:0] ? $signed(coeffs_87) : $signed(_GEN_286);
  wire [31:0] _GEN_288 = 8'h58 == rs2[7:0] ? $signed(coeffs_88) : $signed(_GEN_287);
  wire [31:0] _GEN_289 = 8'h59 == rs2[7:0] ? $signed(coeffs_89) : $signed(_GEN_288);
  wire [31:0] _GEN_290 = 8'h5a == rs2[7:0] ? $signed(coeffs_90) : $signed(_GEN_289);
  wire [31:0] _GEN_291 = 8'h5b == rs2[7:0] ? $signed(coeffs_91) : $signed(_GEN_290);
  wire [31:0] _GEN_292 = 8'h5c == rs2[7:0] ? $signed(coeffs_92) : $signed(_GEN_291);
  wire [31:0] _GEN_293 = 8'h5d == rs2[7:0] ? $signed(coeffs_93) : $signed(_GEN_292);
  wire [31:0] _GEN_294 = 8'h5e == rs2[7:0] ? $signed(coeffs_94) : $signed(_GEN_293);
  wire [31:0] _GEN_295 = 8'h5f == rs2[7:0] ? $signed(coeffs_95) : $signed(_GEN_294);
  wire [31:0] _GEN_296 = 8'h60 == rs2[7:0] ? $signed(coeffs_96) : $signed(_GEN_295);
  wire [31:0] _GEN_297 = 8'h61 == rs2[7:0] ? $signed(coeffs_97) : $signed(_GEN_296);
  wire [31:0] _GEN_298 = 8'h62 == rs2[7:0] ? $signed(coeffs_98) : $signed(_GEN_297);
  wire [31:0] _GEN_299 = 8'h63 == rs2[7:0] ? $signed(coeffs_99) : $signed(_GEN_298);
  wire [31:0] _GEN_300 = 8'h64 == rs2[7:0] ? $signed(coeffs_100) : $signed(_GEN_299);
  wire [31:0] _GEN_301 = 8'h65 == rs2[7:0] ? $signed(coeffs_101) : $signed(_GEN_300);
  wire [31:0] _GEN_302 = 8'h66 == rs2[7:0] ? $signed(coeffs_102) : $signed(_GEN_301);
  wire [31:0] _GEN_303 = 8'h67 == rs2[7:0] ? $signed(coeffs_103) : $signed(_GEN_302);
  wire [31:0] _GEN_304 = 8'h68 == rs2[7:0] ? $signed(coeffs_104) : $signed(_GEN_303);
  wire [31:0] _GEN_305 = 8'h69 == rs2[7:0] ? $signed(coeffs_105) : $signed(_GEN_304);
  wire [31:0] _GEN_306 = 8'h6a == rs2[7:0] ? $signed(coeffs_106) : $signed(_GEN_305);
  wire [31:0] _GEN_307 = 8'h6b == rs2[7:0] ? $signed(coeffs_107) : $signed(_GEN_306);
  wire [31:0] _GEN_308 = 8'h6c == rs2[7:0] ? $signed(coeffs_108) : $signed(_GEN_307);
  wire [31:0] _GEN_309 = 8'h6d == rs2[7:0] ? $signed(coeffs_109) : $signed(_GEN_308);
  wire [31:0] _GEN_310 = 8'h6e == rs2[7:0] ? $signed(coeffs_110) : $signed(_GEN_309);
  wire [31:0] _GEN_311 = 8'h6f == rs2[7:0] ? $signed(coeffs_111) : $signed(_GEN_310);
  wire [31:0] _GEN_312 = 8'h70 == rs2[7:0] ? $signed(coeffs_112) : $signed(_GEN_311);
  wire [31:0] _GEN_313 = 8'h71 == rs2[7:0] ? $signed(coeffs_113) : $signed(_GEN_312);
  wire [31:0] _GEN_314 = 8'h72 == rs2[7:0] ? $signed(coeffs_114) : $signed(_GEN_313);
  wire [31:0] _GEN_315 = 8'h73 == rs2[7:0] ? $signed(coeffs_115) : $signed(_GEN_314);
  wire [31:0] _GEN_316 = 8'h74 == rs2[7:0] ? $signed(coeffs_116) : $signed(_GEN_315);
  wire [31:0] _GEN_317 = 8'h75 == rs2[7:0] ? $signed(coeffs_117) : $signed(_GEN_316);
  wire [31:0] _GEN_318 = 8'h76 == rs2[7:0] ? $signed(coeffs_118) : $signed(_GEN_317);
  wire [31:0] _GEN_319 = 8'h77 == rs2[7:0] ? $signed(coeffs_119) : $signed(_GEN_318);
  wire [31:0] _GEN_320 = 8'h78 == rs2[7:0] ? $signed(coeffs_120) : $signed(_GEN_319);
  wire [31:0] _GEN_321 = 8'h79 == rs2[7:0] ? $signed(coeffs_121) : $signed(_GEN_320);
  wire [31:0] _GEN_322 = 8'h7a == rs2[7:0] ? $signed(coeffs_122) : $signed(_GEN_321);
  wire [31:0] _GEN_323 = 8'h7b == rs2[7:0] ? $signed(coeffs_123) : $signed(_GEN_322);
  wire [31:0] _GEN_324 = 8'h7c == rs2[7:0] ? $signed(coeffs_124) : $signed(_GEN_323);
  wire [31:0] _GEN_325 = 8'h7d == rs2[7:0] ? $signed(coeffs_125) : $signed(_GEN_324);
  wire [31:0] _GEN_326 = 8'h7e == rs2[7:0] ? $signed(coeffs_126) : $signed(_GEN_325);
  wire [31:0] _GEN_327 = 8'h7f == rs2[7:0] ? $signed(coeffs_127) : $signed(_GEN_326);
  wire [31:0] _GEN_328 = 8'h80 == rs2[7:0] ? $signed(coeffs_128) : $signed(_GEN_327);
  wire [31:0] _GEN_329 = 8'h81 == rs2[7:0] ? $signed(coeffs_129) : $signed(_GEN_328);
  wire [31:0] _GEN_330 = 8'h82 == rs2[7:0] ? $signed(coeffs_130) : $signed(_GEN_329);
  wire [31:0] _GEN_331 = 8'h83 == rs2[7:0] ? $signed(coeffs_131) : $signed(_GEN_330);
  wire [31:0] _GEN_332 = 8'h84 == rs2[7:0] ? $signed(coeffs_132) : $signed(_GEN_331);
  wire [31:0] _GEN_333 = 8'h85 == rs2[7:0] ? $signed(coeffs_133) : $signed(_GEN_332);
  wire [31:0] _GEN_334 = 8'h86 == rs2[7:0] ? $signed(coeffs_134) : $signed(_GEN_333);
  wire [31:0] _GEN_335 = 8'h87 == rs2[7:0] ? $signed(coeffs_135) : $signed(_GEN_334);
  wire [31:0] _GEN_336 = 8'h88 == rs2[7:0] ? $signed(coeffs_136) : $signed(_GEN_335);
  wire [31:0] _GEN_337 = 8'h89 == rs2[7:0] ? $signed(coeffs_137) : $signed(_GEN_336);
  wire [31:0] _GEN_338 = 8'h8a == rs2[7:0] ? $signed(coeffs_138) : $signed(_GEN_337);
  wire [31:0] _GEN_339 = 8'h8b == rs2[7:0] ? $signed(coeffs_139) : $signed(_GEN_338);
  wire [31:0] _GEN_340 = 8'h8c == rs2[7:0] ? $signed(coeffs_140) : $signed(_GEN_339);
  wire [31:0] _GEN_341 = 8'h8d == rs2[7:0] ? $signed(coeffs_141) : $signed(_GEN_340);
  wire [31:0] _GEN_342 = 8'h8e == rs2[7:0] ? $signed(coeffs_142) : $signed(_GEN_341);
  wire [31:0] _GEN_343 = 8'h8f == rs2[7:0] ? $signed(coeffs_143) : $signed(_GEN_342);
  wire [31:0] _GEN_344 = 8'h90 == rs2[7:0] ? $signed(coeffs_144) : $signed(_GEN_343);
  wire [31:0] _GEN_345 = 8'h91 == rs2[7:0] ? $signed(coeffs_145) : $signed(_GEN_344);
  wire [31:0] _GEN_346 = 8'h92 == rs2[7:0] ? $signed(coeffs_146) : $signed(_GEN_345);
  wire [31:0] _GEN_347 = 8'h93 == rs2[7:0] ? $signed(coeffs_147) : $signed(_GEN_346);
  wire [31:0] _GEN_348 = 8'h94 == rs2[7:0] ? $signed(coeffs_148) : $signed(_GEN_347);
  wire [31:0] _GEN_349 = 8'h95 == rs2[7:0] ? $signed(coeffs_149) : $signed(_GEN_348);
  wire [31:0] _GEN_350 = 8'h96 == rs2[7:0] ? $signed(coeffs_150) : $signed(_GEN_349);
  wire [31:0] _GEN_351 = 8'h97 == rs2[7:0] ? $signed(coeffs_151) : $signed(_GEN_350);
  wire [31:0] _GEN_352 = 8'h98 == rs2[7:0] ? $signed(coeffs_152) : $signed(_GEN_351);
  wire [31:0] _GEN_353 = 8'h99 == rs2[7:0] ? $signed(coeffs_153) : $signed(_GEN_352);
  wire [31:0] _GEN_354 = 8'h9a == rs2[7:0] ? $signed(coeffs_154) : $signed(_GEN_353);
  wire [31:0] _GEN_355 = 8'h9b == rs2[7:0] ? $signed(coeffs_155) : $signed(_GEN_354);
  wire [31:0] _GEN_356 = 8'h9c == rs2[7:0] ? $signed(coeffs_156) : $signed(_GEN_355);
  wire [31:0] _GEN_357 = 8'h9d == rs2[7:0] ? $signed(coeffs_157) : $signed(_GEN_356);
  wire [31:0] _GEN_358 = 8'h9e == rs2[7:0] ? $signed(coeffs_158) : $signed(_GEN_357);
  wire [31:0] _GEN_359 = 8'h9f == rs2[7:0] ? $signed(coeffs_159) : $signed(_GEN_358);
  wire [31:0] _GEN_360 = 8'ha0 == rs2[7:0] ? $signed(coeffs_160) : $signed(_GEN_359);
  wire [31:0] _GEN_361 = 8'ha1 == rs2[7:0] ? $signed(coeffs_161) : $signed(_GEN_360);
  wire [31:0] _GEN_362 = 8'ha2 == rs2[7:0] ? $signed(coeffs_162) : $signed(_GEN_361);
  wire [31:0] _GEN_363 = 8'ha3 == rs2[7:0] ? $signed(coeffs_163) : $signed(_GEN_362);
  wire [31:0] _GEN_364 = 8'ha4 == rs2[7:0] ? $signed(coeffs_164) : $signed(_GEN_363);
  wire [31:0] _GEN_365 = 8'ha5 == rs2[7:0] ? $signed(coeffs_165) : $signed(_GEN_364);
  wire [31:0] _GEN_366 = 8'ha6 == rs2[7:0] ? $signed(coeffs_166) : $signed(_GEN_365);
  wire [31:0] _GEN_367 = 8'ha7 == rs2[7:0] ? $signed(coeffs_167) : $signed(_GEN_366);
  wire [31:0] _GEN_368 = 8'ha8 == rs2[7:0] ? $signed(coeffs_168) : $signed(_GEN_367);
  wire [31:0] _GEN_369 = 8'ha9 == rs2[7:0] ? $signed(coeffs_169) : $signed(_GEN_368);
  wire [31:0] _GEN_370 = 8'haa == rs2[7:0] ? $signed(coeffs_170) : $signed(_GEN_369);
  wire [31:0] _GEN_371 = 8'hab == rs2[7:0] ? $signed(coeffs_171) : $signed(_GEN_370);
  wire [31:0] _GEN_372 = 8'hac == rs2[7:0] ? $signed(coeffs_172) : $signed(_GEN_371);
  wire [31:0] _GEN_373 = 8'had == rs2[7:0] ? $signed(coeffs_173) : $signed(_GEN_372);
  wire [31:0] _GEN_374 = 8'hae == rs2[7:0] ? $signed(coeffs_174) : $signed(_GEN_373);
  wire [31:0] _GEN_375 = 8'haf == rs2[7:0] ? $signed(coeffs_175) : $signed(_GEN_374);
  wire [31:0] _GEN_376 = 8'hb0 == rs2[7:0] ? $signed(coeffs_176) : $signed(_GEN_375);
  wire [31:0] _GEN_377 = 8'hb1 == rs2[7:0] ? $signed(coeffs_177) : $signed(_GEN_376);
  wire [31:0] _GEN_378 = 8'hb2 == rs2[7:0] ? $signed(coeffs_178) : $signed(_GEN_377);
  wire [31:0] _GEN_379 = 8'hb3 == rs2[7:0] ? $signed(coeffs_179) : $signed(_GEN_378);
  wire [31:0] _GEN_380 = 8'hb4 == rs2[7:0] ? $signed(coeffs_180) : $signed(_GEN_379);
  wire [31:0] _GEN_381 = 8'hb5 == rs2[7:0] ? $signed(coeffs_181) : $signed(_GEN_380);
  wire [31:0] _GEN_382 = 8'hb6 == rs2[7:0] ? $signed(coeffs_182) : $signed(_GEN_381);
  wire [31:0] _GEN_383 = 8'hb7 == rs2[7:0] ? $signed(coeffs_183) : $signed(_GEN_382);
  wire [31:0] _GEN_384 = 8'hb8 == rs2[7:0] ? $signed(coeffs_184) : $signed(_GEN_383);
  wire [31:0] _GEN_385 = 8'hb9 == rs2[7:0] ? $signed(coeffs_185) : $signed(_GEN_384);
  wire [31:0] _GEN_386 = 8'hba == rs2[7:0] ? $signed(coeffs_186) : $signed(_GEN_385);
  wire [31:0] _GEN_387 = 8'hbb == rs2[7:0] ? $signed(coeffs_187) : $signed(_GEN_386);
  wire [31:0] _GEN_388 = 8'hbc == rs2[7:0] ? $signed(coeffs_188) : $signed(_GEN_387);
  wire [31:0] _GEN_389 = 8'hbd == rs2[7:0] ? $signed(coeffs_189) : $signed(_GEN_388);
  wire [31:0] _GEN_390 = 8'hbe == rs2[7:0] ? $signed(coeffs_190) : $signed(_GEN_389);
  wire [31:0] _GEN_391 = 8'hbf == rs2[7:0] ? $signed(coeffs_191) : $signed(_GEN_390);
  wire [31:0] _GEN_392 = 8'hc0 == rs2[7:0] ? $signed(coeffs_192) : $signed(_GEN_391);
  wire [31:0] _GEN_393 = 8'hc1 == rs2[7:0] ? $signed(coeffs_193) : $signed(_GEN_392);
  wire [31:0] _GEN_394 = 8'hc2 == rs2[7:0] ? $signed(coeffs_194) : $signed(_GEN_393);
  wire [31:0] _GEN_395 = 8'hc3 == rs2[7:0] ? $signed(coeffs_195) : $signed(_GEN_394);
  wire [31:0] _GEN_396 = 8'hc4 == rs2[7:0] ? $signed(coeffs_196) : $signed(_GEN_395);
  wire [31:0] _GEN_397 = 8'hc5 == rs2[7:0] ? $signed(coeffs_197) : $signed(_GEN_396);
  wire [31:0] _GEN_398 = 8'hc6 == rs2[7:0] ? $signed(coeffs_198) : $signed(_GEN_397);
  wire [31:0] _GEN_399 = 8'hc7 == rs2[7:0] ? $signed(coeffs_199) : $signed(_GEN_398);
  wire [63:0] _result_T_2 = $signed(data_0) * $signed(coeffs_0);
  wire [63:0] _result_T_3 = $signed(data_1) * $signed(coeffs_1);
  wire [63:0] _result_T_4 = $signed(data_2) * $signed(coeffs_2);
  wire [63:0] _result_T_5 = $signed(data_3) * $signed(coeffs_3);
  wire [63:0] _result_T_6 = $signed(data_4) * $signed(coeffs_4);
  wire [63:0] _result_T_7 = $signed(data_5) * $signed(coeffs_5);
  wire [63:0] _result_T_8 = $signed(data_6) * $signed(coeffs_6);
  wire [63:0] _result_T_9 = $signed(data_7) * $signed(coeffs_7);
  wire [63:0] _result_T_10 = $signed(data_8) * $signed(coeffs_8);
  wire [63:0] _result_T_11 = $signed(data_9) * $signed(coeffs_9);
  wire [63:0] _result_T_12 = $signed(data_10) * $signed(coeffs_10);
  wire [63:0] _result_T_13 = $signed(data_11) * $signed(coeffs_11);
  wire [63:0] _result_T_14 = $signed(data_12) * $signed(coeffs_12);
  wire [63:0] _result_T_15 = $signed(data_13) * $signed(coeffs_13);
  wire [63:0] _result_T_16 = $signed(data_14) * $signed(coeffs_14);
  wire [63:0] _result_T_17 = $signed(data_15) * $signed(coeffs_15);
  wire [63:0] _result_T_18 = $signed(data_16) * $signed(coeffs_16);
  wire [63:0] _result_T_19 = $signed(data_17) * $signed(coeffs_17);
  wire [63:0] _result_T_20 = $signed(data_18) * $signed(coeffs_18);
  wire [63:0] _result_T_21 = $signed(data_19) * $signed(coeffs_19);
  wire [63:0] _result_T_22 = $signed(data_20) * $signed(coeffs_20);
  wire [63:0] _result_T_23 = $signed(data_21) * $signed(coeffs_21);
  wire [63:0] _result_T_24 = $signed(data_22) * $signed(coeffs_22);
  wire [63:0] _result_T_25 = $signed(data_23) * $signed(coeffs_23);
  wire [63:0] _result_T_26 = $signed(data_24) * $signed(coeffs_24);
  wire [63:0] _result_T_27 = $signed(data_25) * $signed(coeffs_25);
  wire [63:0] _result_T_28 = $signed(data_26) * $signed(coeffs_26);
  wire [63:0] _result_T_29 = $signed(data_27) * $signed(coeffs_27);
  wire [63:0] _result_T_30 = $signed(data_28) * $signed(coeffs_28);
  wire [63:0] _result_T_31 = $signed(data_29) * $signed(coeffs_29);
  wire [63:0] _result_T_32 = $signed(data_30) * $signed(coeffs_30);
  wire [63:0] _result_T_33 = $signed(data_31) * $signed(coeffs_31);
  wire [63:0] _result_T_34 = $signed(data_32) * $signed(coeffs_32);
  wire [63:0] _result_T_35 = $signed(data_33) * $signed(coeffs_33);
  wire [63:0] _result_T_36 = $signed(data_34) * $signed(coeffs_34);
  wire [63:0] _result_T_37 = $signed(data_35) * $signed(coeffs_35);
  wire [63:0] _result_T_38 = $signed(data_36) * $signed(coeffs_36);
  wire [63:0] _result_T_39 = $signed(data_37) * $signed(coeffs_37);
  wire [63:0] _result_T_40 = $signed(data_38) * $signed(coeffs_38);
  wire [63:0] _result_T_41 = $signed(data_39) * $signed(coeffs_39);
  wire [63:0] _result_T_42 = $signed(data_40) * $signed(coeffs_40);
  wire [63:0] _result_T_43 = $signed(data_41) * $signed(coeffs_41);
  wire [63:0] _result_T_44 = $signed(data_42) * $signed(coeffs_42);
  wire [63:0] _result_T_45 = $signed(data_43) * $signed(coeffs_43);
  wire [63:0] _result_T_46 = $signed(data_44) * $signed(coeffs_44);
  wire [63:0] _result_T_47 = $signed(data_45) * $signed(coeffs_45);
  wire [63:0] _result_T_48 = $signed(data_46) * $signed(coeffs_46);
  wire [63:0] _result_T_49 = $signed(data_47) * $signed(coeffs_47);
  wire [63:0] _result_T_50 = $signed(data_48) * $signed(coeffs_48);
  wire [63:0] _result_T_51 = $signed(data_49) * $signed(coeffs_49);
  wire [63:0] _result_T_52 = $signed(data_50) * $signed(coeffs_50);
  wire [63:0] _result_T_53 = $signed(data_51) * $signed(coeffs_51);
  wire [63:0] _result_T_54 = $signed(data_52) * $signed(coeffs_52);
  wire [63:0] _result_T_55 = $signed(data_53) * $signed(coeffs_53);
  wire [63:0] _result_T_56 = $signed(data_54) * $signed(coeffs_54);
  wire [63:0] _result_T_57 = $signed(data_55) * $signed(coeffs_55);
  wire [63:0] _result_T_58 = $signed(data_56) * $signed(coeffs_56);
  wire [63:0] _result_T_59 = $signed(data_57) * $signed(coeffs_57);
  wire [63:0] _result_T_60 = $signed(data_58) * $signed(coeffs_58);
  wire [63:0] _result_T_61 = $signed(data_59) * $signed(coeffs_59);
  wire [63:0] _result_T_62 = $signed(data_60) * $signed(coeffs_60);
  wire [63:0] _result_T_63 = $signed(data_61) * $signed(coeffs_61);
  wire [63:0] _result_T_64 = $signed(data_62) * $signed(coeffs_62);
  wire [63:0] _result_T_65 = $signed(data_63) * $signed(coeffs_63);
  wire [63:0] _result_T_66 = $signed(data_64) * $signed(coeffs_64);
  wire [63:0] _result_T_67 = $signed(data_65) * $signed(coeffs_65);
  wire [63:0] _result_T_68 = $signed(data_66) * $signed(coeffs_66);
  wire [63:0] _result_T_69 = $signed(data_67) * $signed(coeffs_67);
  wire [63:0] _result_T_70 = $signed(data_68) * $signed(coeffs_68);
  wire [63:0] _result_T_71 = $signed(data_69) * $signed(coeffs_69);
  wire [63:0] _result_T_72 = $signed(data_70) * $signed(coeffs_70);
  wire [63:0] _result_T_73 = $signed(data_71) * $signed(coeffs_71);
  wire [63:0] _result_T_74 = $signed(data_72) * $signed(coeffs_72);
  wire [63:0] _result_T_75 = $signed(data_73) * $signed(coeffs_73);
  wire [63:0] _result_T_76 = $signed(data_74) * $signed(coeffs_74);
  wire [63:0] _result_T_77 = $signed(data_75) * $signed(coeffs_75);
  wire [63:0] _result_T_78 = $signed(data_76) * $signed(coeffs_76);
  wire [63:0] _result_T_79 = $signed(data_77) * $signed(coeffs_77);
  wire [63:0] _result_T_80 = $signed(data_78) * $signed(coeffs_78);
  wire [63:0] _result_T_81 = $signed(data_79) * $signed(coeffs_79);
  wire [63:0] _result_T_82 = $signed(data_80) * $signed(coeffs_80);
  wire [63:0] _result_T_83 = $signed(data_81) * $signed(coeffs_81);
  wire [63:0] _result_T_84 = $signed(data_82) * $signed(coeffs_82);
  wire [63:0] _result_T_85 = $signed(data_83) * $signed(coeffs_83);
  wire [63:0] _result_T_86 = $signed(data_84) * $signed(coeffs_84);
  wire [63:0] _result_T_87 = $signed(data_85) * $signed(coeffs_85);
  wire [63:0] _result_T_88 = $signed(data_86) * $signed(coeffs_86);
  wire [63:0] _result_T_89 = $signed(data_87) * $signed(coeffs_87);
  wire [63:0] _result_T_90 = $signed(data_88) * $signed(coeffs_88);
  wire [63:0] _result_T_91 = $signed(data_89) * $signed(coeffs_89);
  wire [63:0] _result_T_92 = $signed(data_90) * $signed(coeffs_90);
  wire [63:0] _result_T_93 = $signed(data_91) * $signed(coeffs_91);
  wire [63:0] _result_T_94 = $signed(data_92) * $signed(coeffs_92);
  wire [63:0] _result_T_95 = $signed(data_93) * $signed(coeffs_93);
  wire [63:0] _result_T_96 = $signed(data_94) * $signed(coeffs_94);
  wire [63:0] _result_T_97 = $signed(data_95) * $signed(coeffs_95);
  wire [63:0] _result_T_98 = $signed(data_96) * $signed(coeffs_96);
  wire [63:0] _result_T_99 = $signed(data_97) * $signed(coeffs_97);
  wire [63:0] _result_T_100 = $signed(data_98) * $signed(coeffs_98);
  wire [63:0] _result_T_101 = $signed(data_99) * $signed(coeffs_99);
  wire [63:0] _result_T_102 = $signed(data_100) * $signed(coeffs_100);
  wire [63:0] _result_T_103 = $signed(data_101) * $signed(coeffs_101);
  wire [63:0] _result_T_104 = $signed(data_102) * $signed(coeffs_102);
  wire [63:0] _result_T_105 = $signed(data_103) * $signed(coeffs_103);
  wire [63:0] _result_T_106 = $signed(data_104) * $signed(coeffs_104);
  wire [63:0] _result_T_107 = $signed(data_105) * $signed(coeffs_105);
  wire [63:0] _result_T_108 = $signed(data_106) * $signed(coeffs_106);
  wire [63:0] _result_T_109 = $signed(data_107) * $signed(coeffs_107);
  wire [63:0] _result_T_110 = $signed(data_108) * $signed(coeffs_108);
  wire [63:0] _result_T_111 = $signed(data_109) * $signed(coeffs_109);
  wire [63:0] _result_T_112 = $signed(data_110) * $signed(coeffs_110);
  wire [63:0] _result_T_113 = $signed(data_111) * $signed(coeffs_111);
  wire [63:0] _result_T_114 = $signed(data_112) * $signed(coeffs_112);
  wire [63:0] _result_T_115 = $signed(data_113) * $signed(coeffs_113);
  wire [63:0] _result_T_116 = $signed(data_114) * $signed(coeffs_114);
  wire [63:0] _result_T_117 = $signed(data_115) * $signed(coeffs_115);
  wire [63:0] _result_T_118 = $signed(data_116) * $signed(coeffs_116);
  wire [63:0] _result_T_119 = $signed(data_117) * $signed(coeffs_117);
  wire [63:0] _result_T_120 = $signed(data_118) * $signed(coeffs_118);
  wire [63:0] _result_T_121 = $signed(data_119) * $signed(coeffs_119);
  wire [63:0] _result_T_122 = $signed(data_120) * $signed(coeffs_120);
  wire [63:0] _result_T_123 = $signed(data_121) * $signed(coeffs_121);
  wire [63:0] _result_T_124 = $signed(data_122) * $signed(coeffs_122);
  wire [63:0] _result_T_125 = $signed(data_123) * $signed(coeffs_123);
  wire [63:0] _result_T_126 = $signed(data_124) * $signed(coeffs_124);
  wire [63:0] _result_T_127 = $signed(data_125) * $signed(coeffs_125);
  wire [63:0] _result_T_128 = $signed(data_126) * $signed(coeffs_126);
  wire [63:0] _result_T_129 = $signed(data_127) * $signed(coeffs_127);
  wire [63:0] _result_T_130 = $signed(data_128) * $signed(coeffs_128);
  wire [63:0] _result_T_131 = $signed(data_129) * $signed(coeffs_129);
  wire [63:0] _result_T_132 = $signed(data_130) * $signed(coeffs_130);
  wire [63:0] _result_T_133 = $signed(data_131) * $signed(coeffs_131);
  wire [63:0] _result_T_134 = $signed(data_132) * $signed(coeffs_132);
  wire [63:0] _result_T_135 = $signed(data_133) * $signed(coeffs_133);
  wire [63:0] _result_T_136 = $signed(data_134) * $signed(coeffs_134);
  wire [63:0] _result_T_137 = $signed(data_135) * $signed(coeffs_135);
  wire [63:0] _result_T_138 = $signed(data_136) * $signed(coeffs_136);
  wire [63:0] _result_T_139 = $signed(data_137) * $signed(coeffs_137);
  wire [63:0] _result_T_140 = $signed(data_138) * $signed(coeffs_138);
  wire [63:0] _result_T_141 = $signed(data_139) * $signed(coeffs_139);
  wire [63:0] _result_T_142 = $signed(data_140) * $signed(coeffs_140);
  wire [63:0] _result_T_143 = $signed(data_141) * $signed(coeffs_141);
  wire [63:0] _result_T_144 = $signed(data_142) * $signed(coeffs_142);
  wire [63:0] _result_T_145 = $signed(data_143) * $signed(coeffs_143);
  wire [63:0] _result_T_146 = $signed(data_144) * $signed(coeffs_144);
  wire [63:0] _result_T_147 = $signed(data_145) * $signed(coeffs_145);
  wire [63:0] _result_T_148 = $signed(data_146) * $signed(coeffs_146);
  wire [63:0] _result_T_149 = $signed(data_147) * $signed(coeffs_147);
  wire [63:0] _result_T_150 = $signed(data_148) * $signed(coeffs_148);
  wire [63:0] _result_T_151 = $signed(data_149) * $signed(coeffs_149);
  wire [63:0] _result_T_152 = $signed(data_150) * $signed(coeffs_150);
  wire [63:0] _result_T_153 = $signed(data_151) * $signed(coeffs_151);
  wire [63:0] _result_T_154 = $signed(data_152) * $signed(coeffs_152);
  wire [63:0] _result_T_155 = $signed(data_153) * $signed(coeffs_153);
  wire [63:0] _result_T_156 = $signed(data_154) * $signed(coeffs_154);
  wire [63:0] _result_T_157 = $signed(data_155) * $signed(coeffs_155);
  wire [63:0] _result_T_158 = $signed(data_156) * $signed(coeffs_156);
  wire [63:0] _result_T_159 = $signed(data_157) * $signed(coeffs_157);
  wire [63:0] _result_T_160 = $signed(data_158) * $signed(coeffs_158);
  wire [63:0] _result_T_161 = $signed(data_159) * $signed(coeffs_159);
  wire [63:0] _result_T_162 = $signed(data_160) * $signed(coeffs_160);
  wire [63:0] _result_T_163 = $signed(data_161) * $signed(coeffs_161);
  wire [63:0] _result_T_164 = $signed(data_162) * $signed(coeffs_162);
  wire [63:0] _result_T_165 = $signed(data_163) * $signed(coeffs_163);
  wire [63:0] _result_T_166 = $signed(data_164) * $signed(coeffs_164);
  wire [63:0] _result_T_167 = $signed(data_165) * $signed(coeffs_165);
  wire [63:0] _result_T_168 = $signed(data_166) * $signed(coeffs_166);
  wire [63:0] _result_T_169 = $signed(data_167) * $signed(coeffs_167);
  wire [63:0] _result_T_170 = $signed(data_168) * $signed(coeffs_168);
  wire [63:0] _result_T_171 = $signed(data_169) * $signed(coeffs_169);
  wire [63:0] _result_T_172 = $signed(data_170) * $signed(coeffs_170);
  wire [63:0] _result_T_173 = $signed(data_171) * $signed(coeffs_171);
  wire [63:0] _result_T_174 = $signed(data_172) * $signed(coeffs_172);
  wire [63:0] _result_T_175 = $signed(data_173) * $signed(coeffs_173);
  wire [63:0] _result_T_176 = $signed(data_174) * $signed(coeffs_174);
  wire [63:0] _result_T_177 = $signed(data_175) * $signed(coeffs_175);
  wire [63:0] _result_T_178 = $signed(data_176) * $signed(coeffs_176);
  wire [63:0] _result_T_179 = $signed(data_177) * $signed(coeffs_177);
  wire [63:0] _result_T_180 = $signed(data_178) * $signed(coeffs_178);
  wire [63:0] _result_T_181 = $signed(data_179) * $signed(coeffs_179);
  wire [63:0] _result_T_182 = $signed(data_180) * $signed(coeffs_180);
  wire [63:0] _result_T_183 = $signed(data_181) * $signed(coeffs_181);
  wire [63:0] _result_T_184 = $signed(data_182) * $signed(coeffs_182);
  wire [63:0] _result_T_185 = $signed(data_183) * $signed(coeffs_183);
  wire [63:0] _result_T_186 = $signed(data_184) * $signed(coeffs_184);
  wire [63:0] _result_T_187 = $signed(data_185) * $signed(coeffs_185);
  wire [63:0] _result_T_188 = $signed(data_186) * $signed(coeffs_186);
  wire [63:0] _result_T_189 = $signed(data_187) * $signed(coeffs_187);
  wire [63:0] _result_T_190 = $signed(data_188) * $signed(coeffs_188);
  wire [63:0] _result_T_191 = $signed(data_189) * $signed(coeffs_189);
  wire [63:0] _result_T_192 = $signed(data_190) * $signed(coeffs_190);
  wire [63:0] _result_T_193 = $signed(data_191) * $signed(coeffs_191);
  wire [63:0] _result_T_194 = $signed(data_192) * $signed(coeffs_192);
  wire [63:0] _result_T_195 = $signed(data_193) * $signed(coeffs_193);
  wire [63:0] _result_T_196 = $signed(data_194) * $signed(coeffs_194);
  wire [63:0] _result_T_197 = $signed(data_195) * $signed(coeffs_195);
  wire [63:0] _result_T_198 = $signed(data_196) * $signed(coeffs_196);
  wire [63:0] _result_T_199 = $signed(data_197) * $signed(coeffs_197);
  wire [63:0] _result_T_200 = $signed(data_198) * $signed(coeffs_198);
  wire [63:0] _result_T_201 = $signed(data_199) * $signed(coeffs_199);
  wire [63:0] _result_T_204 = $signed(_result_T_2) + $signed(_result_T_3);
  wire [63:0] _result_T_207 = $signed(_result_T_204) + $signed(_result_T_4);
  wire [63:0] _result_T_210 = $signed(_result_T_207) + $signed(_result_T_5);
  wire [63:0] _result_T_213 = $signed(_result_T_210) + $signed(_result_T_6);
  wire [63:0] _result_T_216 = $signed(_result_T_213) + $signed(_result_T_7);
  wire [63:0] _result_T_219 = $signed(_result_T_216) + $signed(_result_T_8);
  wire [63:0] _result_T_222 = $signed(_result_T_219) + $signed(_result_T_9);
  wire [63:0] _result_T_225 = $signed(_result_T_222) + $signed(_result_T_10);
  wire [63:0] _result_T_228 = $signed(_result_T_225) + $signed(_result_T_11);
  wire [63:0] _result_T_231 = $signed(_result_T_228) + $signed(_result_T_12);
  wire [63:0] _result_T_234 = $signed(_result_T_231) + $signed(_result_T_13);
  wire [63:0] _result_T_237 = $signed(_result_T_234) + $signed(_result_T_14);
  wire [63:0] _result_T_240 = $signed(_result_T_237) + $signed(_result_T_15);
  wire [63:0] _result_T_243 = $signed(_result_T_240) + $signed(_result_T_16);
  wire [63:0] _result_T_246 = $signed(_result_T_243) + $signed(_result_T_17);
  wire [63:0] _result_T_249 = $signed(_result_T_246) + $signed(_result_T_18);
  wire [63:0] _result_T_252 = $signed(_result_T_249) + $signed(_result_T_19);
  wire [63:0] _result_T_255 = $signed(_result_T_252) + $signed(_result_T_20);
  wire [63:0] _result_T_258 = $signed(_result_T_255) + $signed(_result_T_21);
  wire [63:0] _result_T_261 = $signed(_result_T_258) + $signed(_result_T_22);
  wire [63:0] _result_T_264 = $signed(_result_T_261) + $signed(_result_T_23);
  wire [63:0] _result_T_267 = $signed(_result_T_264) + $signed(_result_T_24);
  wire [63:0] _result_T_270 = $signed(_result_T_267) + $signed(_result_T_25);
  wire [63:0] _result_T_273 = $signed(_result_T_270) + $signed(_result_T_26);
  wire [63:0] _result_T_276 = $signed(_result_T_273) + $signed(_result_T_27);
  wire [63:0] _result_T_279 = $signed(_result_T_276) + $signed(_result_T_28);
  wire [63:0] _result_T_282 = $signed(_result_T_279) + $signed(_result_T_29);
  wire [63:0] _result_T_285 = $signed(_result_T_282) + $signed(_result_T_30);
  wire [63:0] _result_T_288 = $signed(_result_T_285) + $signed(_result_T_31);
  wire [63:0] _result_T_291 = $signed(_result_T_288) + $signed(_result_T_32);
  wire [63:0] _result_T_294 = $signed(_result_T_291) + $signed(_result_T_33);
  wire [63:0] _result_T_297 = $signed(_result_T_294) + $signed(_result_T_34);
  wire [63:0] _result_T_300 = $signed(_result_T_297) + $signed(_result_T_35);
  wire [63:0] _result_T_303 = $signed(_result_T_300) + $signed(_result_T_36);
  wire [63:0] _result_T_306 = $signed(_result_T_303) + $signed(_result_T_37);
  wire [63:0] _result_T_309 = $signed(_result_T_306) + $signed(_result_T_38);
  wire [63:0] _result_T_312 = $signed(_result_T_309) + $signed(_result_T_39);
  wire [63:0] _result_T_315 = $signed(_result_T_312) + $signed(_result_T_40);
  wire [63:0] _result_T_318 = $signed(_result_T_315) + $signed(_result_T_41);
  wire [63:0] _result_T_321 = $signed(_result_T_318) + $signed(_result_T_42);
  wire [63:0] _result_T_324 = $signed(_result_T_321) + $signed(_result_T_43);
  wire [63:0] _result_T_327 = $signed(_result_T_324) + $signed(_result_T_44);
  wire [63:0] _result_T_330 = $signed(_result_T_327) + $signed(_result_T_45);
  wire [63:0] _result_T_333 = $signed(_result_T_330) + $signed(_result_T_46);
  wire [63:0] _result_T_336 = $signed(_result_T_333) + $signed(_result_T_47);
  wire [63:0] _result_T_339 = $signed(_result_T_336) + $signed(_result_T_48);
  wire [63:0] _result_T_342 = $signed(_result_T_339) + $signed(_result_T_49);
  wire [63:0] _result_T_345 = $signed(_result_T_342) + $signed(_result_T_50);
  wire [63:0] _result_T_348 = $signed(_result_T_345) + $signed(_result_T_51);
  wire [63:0] _result_T_351 = $signed(_result_T_348) + $signed(_result_T_52);
  wire [63:0] _result_T_354 = $signed(_result_T_351) + $signed(_result_T_53);
  wire [63:0] _result_T_357 = $signed(_result_T_354) + $signed(_result_T_54);
  wire [63:0] _result_T_360 = $signed(_result_T_357) + $signed(_result_T_55);
  wire [63:0] _result_T_363 = $signed(_result_T_360) + $signed(_result_T_56);
  wire [63:0] _result_T_366 = $signed(_result_T_363) + $signed(_result_T_57);
  wire [63:0] _result_T_369 = $signed(_result_T_366) + $signed(_result_T_58);
  wire [63:0] _result_T_372 = $signed(_result_T_369) + $signed(_result_T_59);
  wire [63:0] _result_T_375 = $signed(_result_T_372) + $signed(_result_T_60);
  wire [63:0] _result_T_378 = $signed(_result_T_375) + $signed(_result_T_61);
  wire [63:0] _result_T_381 = $signed(_result_T_378) + $signed(_result_T_62);
  wire [63:0] _result_T_384 = $signed(_result_T_381) + $signed(_result_T_63);
  wire [63:0] _result_T_387 = $signed(_result_T_384) + $signed(_result_T_64);
  wire [63:0] _result_T_390 = $signed(_result_T_387) + $signed(_result_T_65);
  wire [63:0] _result_T_393 = $signed(_result_T_390) + $signed(_result_T_66);
  wire [63:0] _result_T_396 = $signed(_result_T_393) + $signed(_result_T_67);
  wire [63:0] _result_T_399 = $signed(_result_T_396) + $signed(_result_T_68);
  wire [63:0] _result_T_402 = $signed(_result_T_399) + $signed(_result_T_69);
  wire [63:0] _result_T_405 = $signed(_result_T_402) + $signed(_result_T_70);
  wire [63:0] _result_T_408 = $signed(_result_T_405) + $signed(_result_T_71);
  wire [63:0] _result_T_411 = $signed(_result_T_408) + $signed(_result_T_72);
  wire [63:0] _result_T_414 = $signed(_result_T_411) + $signed(_result_T_73);
  wire [63:0] _result_T_417 = $signed(_result_T_414) + $signed(_result_T_74);
  wire [63:0] _result_T_420 = $signed(_result_T_417) + $signed(_result_T_75);
  wire [63:0] _result_T_423 = $signed(_result_T_420) + $signed(_result_T_76);
  wire [63:0] _result_T_426 = $signed(_result_T_423) + $signed(_result_T_77);
  wire [63:0] _result_T_429 = $signed(_result_T_426) + $signed(_result_T_78);
  wire [63:0] _result_T_432 = $signed(_result_T_429) + $signed(_result_T_79);
  wire [63:0] _result_T_435 = $signed(_result_T_432) + $signed(_result_T_80);
  wire [63:0] _result_T_438 = $signed(_result_T_435) + $signed(_result_T_81);
  wire [63:0] _result_T_441 = $signed(_result_T_438) + $signed(_result_T_82);
  wire [63:0] _result_T_444 = $signed(_result_T_441) + $signed(_result_T_83);
  wire [63:0] _result_T_447 = $signed(_result_T_444) + $signed(_result_T_84);
  wire [63:0] _result_T_450 = $signed(_result_T_447) + $signed(_result_T_85);
  wire [63:0] _result_T_453 = $signed(_result_T_450) + $signed(_result_T_86);
  wire [63:0] _result_T_456 = $signed(_result_T_453) + $signed(_result_T_87);
  wire [63:0] _result_T_459 = $signed(_result_T_456) + $signed(_result_T_88);
  wire [63:0] _result_T_462 = $signed(_result_T_459) + $signed(_result_T_89);
  wire [63:0] _result_T_465 = $signed(_result_T_462) + $signed(_result_T_90);
  wire [63:0] _result_T_468 = $signed(_result_T_465) + $signed(_result_T_91);
  wire [63:0] _result_T_471 = $signed(_result_T_468) + $signed(_result_T_92);
  wire [63:0] _result_T_474 = $signed(_result_T_471) + $signed(_result_T_93);
  wire [63:0] _result_T_477 = $signed(_result_T_474) + $signed(_result_T_94);
  wire [63:0] _result_T_480 = $signed(_result_T_477) + $signed(_result_T_95);
  wire [63:0] _result_T_483 = $signed(_result_T_480) + $signed(_result_T_96);
  wire [63:0] _result_T_486 = $signed(_result_T_483) + $signed(_result_T_97);
  wire [63:0] _result_T_489 = $signed(_result_T_486) + $signed(_result_T_98);
  wire [63:0] _result_T_492 = $signed(_result_T_489) + $signed(_result_T_99);
  wire [63:0] _result_T_495 = $signed(_result_T_492) + $signed(_result_T_100);
  wire [63:0] _result_T_498 = $signed(_result_T_495) + $signed(_result_T_101);
  wire [63:0] _result_T_501 = $signed(_result_T_498) + $signed(_result_T_102);
  wire [63:0] _result_T_504 = $signed(_result_T_501) + $signed(_result_T_103);
  wire [63:0] _result_T_507 = $signed(_result_T_504) + $signed(_result_T_104);
  wire [63:0] _result_T_510 = $signed(_result_T_507) + $signed(_result_T_105);
  wire [63:0] _result_T_513 = $signed(_result_T_510) + $signed(_result_T_106);
  wire [63:0] _result_T_516 = $signed(_result_T_513) + $signed(_result_T_107);
  wire [63:0] _result_T_519 = $signed(_result_T_516) + $signed(_result_T_108);
  wire [63:0] _result_T_522 = $signed(_result_T_519) + $signed(_result_T_109);
  wire [63:0] _result_T_525 = $signed(_result_T_522) + $signed(_result_T_110);
  wire [63:0] _result_T_528 = $signed(_result_T_525) + $signed(_result_T_111);
  wire [63:0] _result_T_531 = $signed(_result_T_528) + $signed(_result_T_112);
  wire [63:0] _result_T_534 = $signed(_result_T_531) + $signed(_result_T_113);
  wire [63:0] _result_T_537 = $signed(_result_T_534) + $signed(_result_T_114);
  wire [63:0] _result_T_540 = $signed(_result_T_537) + $signed(_result_T_115);
  wire [63:0] _result_T_543 = $signed(_result_T_540) + $signed(_result_T_116);
  wire [63:0] _result_T_546 = $signed(_result_T_543) + $signed(_result_T_117);
  wire [63:0] _result_T_549 = $signed(_result_T_546) + $signed(_result_T_118);
  wire [63:0] _result_T_552 = $signed(_result_T_549) + $signed(_result_T_119);
  wire [63:0] _result_T_555 = $signed(_result_T_552) + $signed(_result_T_120);
  wire [63:0] _result_T_558 = $signed(_result_T_555) + $signed(_result_T_121);
  wire [63:0] _result_T_561 = $signed(_result_T_558) + $signed(_result_T_122);
  wire [63:0] _result_T_564 = $signed(_result_T_561) + $signed(_result_T_123);
  wire [63:0] _result_T_567 = $signed(_result_T_564) + $signed(_result_T_124);
  wire [63:0] _result_T_570 = $signed(_result_T_567) + $signed(_result_T_125);
  wire [63:0] _result_T_573 = $signed(_result_T_570) + $signed(_result_T_126);
  wire [63:0] _result_T_576 = $signed(_result_T_573) + $signed(_result_T_127);
  wire [63:0] _result_T_579 = $signed(_result_T_576) + $signed(_result_T_128);
  wire [63:0] _result_T_582 = $signed(_result_T_579) + $signed(_result_T_129);
  wire [63:0] _result_T_585 = $signed(_result_T_582) + $signed(_result_T_130);
  wire [63:0] _result_T_588 = $signed(_result_T_585) + $signed(_result_T_131);
  wire [63:0] _result_T_591 = $signed(_result_T_588) + $signed(_result_T_132);
  wire [63:0] _result_T_594 = $signed(_result_T_591) + $signed(_result_T_133);
  wire [63:0] _result_T_597 = $signed(_result_T_594) + $signed(_result_T_134);
  wire [63:0] _result_T_600 = $signed(_result_T_597) + $signed(_result_T_135);
  wire [63:0] _result_T_603 = $signed(_result_T_600) + $signed(_result_T_136);
  wire [63:0] _result_T_606 = $signed(_result_T_603) + $signed(_result_T_137);
  wire [63:0] _result_T_609 = $signed(_result_T_606) + $signed(_result_T_138);
  wire [63:0] _result_T_612 = $signed(_result_T_609) + $signed(_result_T_139);
  wire [63:0] _result_T_615 = $signed(_result_T_612) + $signed(_result_T_140);
  wire [63:0] _result_T_618 = $signed(_result_T_615) + $signed(_result_T_141);
  wire [63:0] _result_T_621 = $signed(_result_T_618) + $signed(_result_T_142);
  wire [63:0] _result_T_624 = $signed(_result_T_621) + $signed(_result_T_143);
  wire [63:0] _result_T_627 = $signed(_result_T_624) + $signed(_result_T_144);
  wire [63:0] _result_T_630 = $signed(_result_T_627) + $signed(_result_T_145);
  wire [63:0] _result_T_633 = $signed(_result_T_630) + $signed(_result_T_146);
  wire [63:0] _result_T_636 = $signed(_result_T_633) + $signed(_result_T_147);
  wire [63:0] _result_T_639 = $signed(_result_T_636) + $signed(_result_T_148);
  wire [63:0] _result_T_642 = $signed(_result_T_639) + $signed(_result_T_149);
  wire [63:0] _result_T_645 = $signed(_result_T_642) + $signed(_result_T_150);
  wire [63:0] _result_T_648 = $signed(_result_T_645) + $signed(_result_T_151);
  wire [63:0] _result_T_651 = $signed(_result_T_648) + $signed(_result_T_152);
  wire [63:0] _result_T_654 = $signed(_result_T_651) + $signed(_result_T_153);
  wire [63:0] _result_T_657 = $signed(_result_T_654) + $signed(_result_T_154);
  wire [63:0] _result_T_660 = $signed(_result_T_657) + $signed(_result_T_155);
  wire [63:0] _result_T_663 = $signed(_result_T_660) + $signed(_result_T_156);
  wire [63:0] _result_T_666 = $signed(_result_T_663) + $signed(_result_T_157);
  wire [63:0] _result_T_669 = $signed(_result_T_666) + $signed(_result_T_158);
  wire [63:0] _result_T_672 = $signed(_result_T_669) + $signed(_result_T_159);
  wire [63:0] _result_T_675 = $signed(_result_T_672) + $signed(_result_T_160);
  wire [63:0] _result_T_678 = $signed(_result_T_675) + $signed(_result_T_161);
  wire [63:0] _result_T_681 = $signed(_result_T_678) + $signed(_result_T_162);
  wire [63:0] _result_T_684 = $signed(_result_T_681) + $signed(_result_T_163);
  wire [63:0] _result_T_687 = $signed(_result_T_684) + $signed(_result_T_164);
  wire [63:0] _result_T_690 = $signed(_result_T_687) + $signed(_result_T_165);
  wire [63:0] _result_T_693 = $signed(_result_T_690) + $signed(_result_T_166);
  wire [63:0] _result_T_696 = $signed(_result_T_693) + $signed(_result_T_167);
  wire [63:0] _result_T_699 = $signed(_result_T_696) + $signed(_result_T_168);
  wire [63:0] _result_T_702 = $signed(_result_T_699) + $signed(_result_T_169);
  wire [63:0] _result_T_705 = $signed(_result_T_702) + $signed(_result_T_170);
  wire [63:0] _result_T_708 = $signed(_result_T_705) + $signed(_result_T_171);
  wire [63:0] _result_T_711 = $signed(_result_T_708) + $signed(_result_T_172);
  wire [63:0] _result_T_714 = $signed(_result_T_711) + $signed(_result_T_173);
  wire [63:0] _result_T_717 = $signed(_result_T_714) + $signed(_result_T_174);
  wire [63:0] _result_T_720 = $signed(_result_T_717) + $signed(_result_T_175);
  wire [63:0] _result_T_723 = $signed(_result_T_720) + $signed(_result_T_176);
  wire [63:0] _result_T_726 = $signed(_result_T_723) + $signed(_result_T_177);
  wire [63:0] _result_T_729 = $signed(_result_T_726) + $signed(_result_T_178);
  wire [63:0] _result_T_732 = $signed(_result_T_729) + $signed(_result_T_179);
  wire [63:0] _result_T_735 = $signed(_result_T_732) + $signed(_result_T_180);
  wire [63:0] _result_T_738 = $signed(_result_T_735) + $signed(_result_T_181);
  wire [63:0] _result_T_741 = $signed(_result_T_738) + $signed(_result_T_182);
  wire [63:0] _result_T_744 = $signed(_result_T_741) + $signed(_result_T_183);
  wire [63:0] _result_T_747 = $signed(_result_T_744) + $signed(_result_T_184);
  wire [63:0] _result_T_750 = $signed(_result_T_747) + $signed(_result_T_185);
  wire [63:0] _result_T_753 = $signed(_result_T_750) + $signed(_result_T_186);
  wire [63:0] _result_T_756 = $signed(_result_T_753) + $signed(_result_T_187);
  wire [63:0] _result_T_759 = $signed(_result_T_756) + $signed(_result_T_188);
  wire [63:0] _result_T_762 = $signed(_result_T_759) + $signed(_result_T_189);
  wire [63:0] _result_T_765 = $signed(_result_T_762) + $signed(_result_T_190);
  wire [63:0] _result_T_768 = $signed(_result_T_765) + $signed(_result_T_191);
  wire [63:0] _result_T_771 = $signed(_result_T_768) + $signed(_result_T_192);
  wire [63:0] _result_T_774 = $signed(_result_T_771) + $signed(_result_T_193);
  wire [63:0] _result_T_777 = $signed(_result_T_774) + $signed(_result_T_194);
  wire [63:0] _result_T_780 = $signed(_result_T_777) + $signed(_result_T_195);
  wire [63:0] _result_T_783 = $signed(_result_T_780) + $signed(_result_T_196);
  wire [63:0] _result_T_786 = $signed(_result_T_783) + $signed(_result_T_197);
  wire [63:0] _result_T_789 = $signed(_result_T_786) + $signed(_result_T_198);
  wire [63:0] _result_T_792 = $signed(_result_T_789) + $signed(_result_T_199);
  wire [63:0] _result_T_795 = $signed(_result_T_792) + $signed(_result_T_200);
  wire [63:0] _result_T_798 = $signed(_result_T_795) + $signed(_result_T_201);
  wire [63:0] _GEN_400 = insn[6:0] == 7'h3b ? $signed(_result_T_798) : $signed(result);
  assign rd = result[31:0];
  always @(posedge clock) begin
    if (reset) begin
      coeffs_0 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h0 == rs2[7:0]) begin
          coeffs_0 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_1 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h1 == rs2[7:0]) begin
          coeffs_1 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_2 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h2 == rs2[7:0]) begin
          coeffs_2 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_3 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h3 == rs2[7:0]) begin
          coeffs_3 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_4 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h4 == rs2[7:0]) begin
          coeffs_4 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_5 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h5 == rs2[7:0]) begin
          coeffs_5 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_6 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h6 == rs2[7:0]) begin
          coeffs_6 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_7 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h7 == rs2[7:0]) begin
          coeffs_7 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_8 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h8 == rs2[7:0]) begin
          coeffs_8 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_9 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h9 == rs2[7:0]) begin
          coeffs_9 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_10 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'ha == rs2[7:0]) begin
          coeffs_10 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_11 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hb == rs2[7:0]) begin
          coeffs_11 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_12 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hc == rs2[7:0]) begin
          coeffs_12 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_13 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hd == rs2[7:0]) begin
          coeffs_13 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_14 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'he == rs2[7:0]) begin
          coeffs_14 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_15 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hf == rs2[7:0]) begin
          coeffs_15 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_16 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h10 == rs2[7:0]) begin
          coeffs_16 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_17 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h11 == rs2[7:0]) begin
          coeffs_17 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_18 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h12 == rs2[7:0]) begin
          coeffs_18 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_19 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h13 == rs2[7:0]) begin
          coeffs_19 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_20 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h14 == rs2[7:0]) begin
          coeffs_20 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_21 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h15 == rs2[7:0]) begin
          coeffs_21 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_22 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h16 == rs2[7:0]) begin
          coeffs_22 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_23 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h17 == rs2[7:0]) begin
          coeffs_23 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_24 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h18 == rs2[7:0]) begin
          coeffs_24 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_25 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h19 == rs2[7:0]) begin
          coeffs_25 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_26 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h1a == rs2[7:0]) begin
          coeffs_26 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_27 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h1b == rs2[7:0]) begin
          coeffs_27 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_28 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h1c == rs2[7:0]) begin
          coeffs_28 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_29 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h1d == rs2[7:0]) begin
          coeffs_29 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_30 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h1e == rs2[7:0]) begin
          coeffs_30 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_31 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h1f == rs2[7:0]) begin
          coeffs_31 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_32 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h20 == rs2[7:0]) begin
          coeffs_32 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_33 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h21 == rs2[7:0]) begin
          coeffs_33 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_34 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h22 == rs2[7:0]) begin
          coeffs_34 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_35 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h23 == rs2[7:0]) begin
          coeffs_35 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_36 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h24 == rs2[7:0]) begin
          coeffs_36 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_37 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h25 == rs2[7:0]) begin
          coeffs_37 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_38 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h26 == rs2[7:0]) begin
          coeffs_38 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_39 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h27 == rs2[7:0]) begin
          coeffs_39 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_40 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h28 == rs2[7:0]) begin
          coeffs_40 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_41 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h29 == rs2[7:0]) begin
          coeffs_41 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_42 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h2a == rs2[7:0]) begin
          coeffs_42 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_43 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h2b == rs2[7:0]) begin
          coeffs_43 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_44 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h2c == rs2[7:0]) begin
          coeffs_44 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_45 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h2d == rs2[7:0]) begin
          coeffs_45 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_46 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h2e == rs2[7:0]) begin
          coeffs_46 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_47 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h2f == rs2[7:0]) begin
          coeffs_47 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_48 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h30 == rs2[7:0]) begin
          coeffs_48 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_49 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h31 == rs2[7:0]) begin
          coeffs_49 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_50 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h32 == rs2[7:0]) begin
          coeffs_50 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_51 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h33 == rs2[7:0]) begin
          coeffs_51 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_52 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h34 == rs2[7:0]) begin
          coeffs_52 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_53 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h35 == rs2[7:0]) begin
          coeffs_53 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_54 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h36 == rs2[7:0]) begin
          coeffs_54 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_55 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h37 == rs2[7:0]) begin
          coeffs_55 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_56 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h38 == rs2[7:0]) begin
          coeffs_56 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_57 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h39 == rs2[7:0]) begin
          coeffs_57 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_58 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h3a == rs2[7:0]) begin
          coeffs_58 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_59 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h3b == rs2[7:0]) begin
          coeffs_59 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_60 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h3c == rs2[7:0]) begin
          coeffs_60 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_61 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h3d == rs2[7:0]) begin
          coeffs_61 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_62 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h3e == rs2[7:0]) begin
          coeffs_62 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_63 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h3f == rs2[7:0]) begin
          coeffs_63 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_64 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h40 == rs2[7:0]) begin
          coeffs_64 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_65 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h41 == rs2[7:0]) begin
          coeffs_65 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_66 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h42 == rs2[7:0]) begin
          coeffs_66 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_67 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h43 == rs2[7:0]) begin
          coeffs_67 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_68 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h44 == rs2[7:0]) begin
          coeffs_68 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_69 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h45 == rs2[7:0]) begin
          coeffs_69 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_70 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h46 == rs2[7:0]) begin
          coeffs_70 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_71 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h47 == rs2[7:0]) begin
          coeffs_71 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_72 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h48 == rs2[7:0]) begin
          coeffs_72 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_73 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h49 == rs2[7:0]) begin
          coeffs_73 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_74 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h4a == rs2[7:0]) begin
          coeffs_74 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_75 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h4b == rs2[7:0]) begin
          coeffs_75 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_76 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h4c == rs2[7:0]) begin
          coeffs_76 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_77 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h4d == rs2[7:0]) begin
          coeffs_77 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_78 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h4e == rs2[7:0]) begin
          coeffs_78 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_79 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h4f == rs2[7:0]) begin
          coeffs_79 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_80 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h50 == rs2[7:0]) begin
          coeffs_80 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_81 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h51 == rs2[7:0]) begin
          coeffs_81 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_82 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h52 == rs2[7:0]) begin
          coeffs_82 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_83 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h53 == rs2[7:0]) begin
          coeffs_83 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_84 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h54 == rs2[7:0]) begin
          coeffs_84 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_85 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h55 == rs2[7:0]) begin
          coeffs_85 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_86 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h56 == rs2[7:0]) begin
          coeffs_86 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_87 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h57 == rs2[7:0]) begin
          coeffs_87 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_88 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h58 == rs2[7:0]) begin
          coeffs_88 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_89 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h59 == rs2[7:0]) begin
          coeffs_89 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_90 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h5a == rs2[7:0]) begin
          coeffs_90 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_91 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h5b == rs2[7:0]) begin
          coeffs_91 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_92 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h5c == rs2[7:0]) begin
          coeffs_92 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_93 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h5d == rs2[7:0]) begin
          coeffs_93 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_94 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h5e == rs2[7:0]) begin
          coeffs_94 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_95 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h5f == rs2[7:0]) begin
          coeffs_95 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_96 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h60 == rs2[7:0]) begin
          coeffs_96 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_97 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h61 == rs2[7:0]) begin
          coeffs_97 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_98 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h62 == rs2[7:0]) begin
          coeffs_98 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_99 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h63 == rs2[7:0]) begin
          coeffs_99 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_100 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h64 == rs2[7:0]) begin
          coeffs_100 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_101 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h65 == rs2[7:0]) begin
          coeffs_101 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_102 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h66 == rs2[7:0]) begin
          coeffs_102 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_103 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h67 == rs2[7:0]) begin
          coeffs_103 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_104 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h68 == rs2[7:0]) begin
          coeffs_104 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_105 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h69 == rs2[7:0]) begin
          coeffs_105 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_106 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h6a == rs2[7:0]) begin
          coeffs_106 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_107 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h6b == rs2[7:0]) begin
          coeffs_107 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_108 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h6c == rs2[7:0]) begin
          coeffs_108 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_109 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h6d == rs2[7:0]) begin
          coeffs_109 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_110 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h6e == rs2[7:0]) begin
          coeffs_110 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_111 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h6f == rs2[7:0]) begin
          coeffs_111 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_112 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h70 == rs2[7:0]) begin
          coeffs_112 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_113 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h71 == rs2[7:0]) begin
          coeffs_113 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_114 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h72 == rs2[7:0]) begin
          coeffs_114 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_115 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h73 == rs2[7:0]) begin
          coeffs_115 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_116 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h74 == rs2[7:0]) begin
          coeffs_116 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_117 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h75 == rs2[7:0]) begin
          coeffs_117 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_118 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h76 == rs2[7:0]) begin
          coeffs_118 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_119 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h77 == rs2[7:0]) begin
          coeffs_119 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_120 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h78 == rs2[7:0]) begin
          coeffs_120 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_121 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h79 == rs2[7:0]) begin
          coeffs_121 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_122 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h7a == rs2[7:0]) begin
          coeffs_122 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_123 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h7b == rs2[7:0]) begin
          coeffs_123 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_124 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h7c == rs2[7:0]) begin
          coeffs_124 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_125 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h7d == rs2[7:0]) begin
          coeffs_125 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_126 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h7e == rs2[7:0]) begin
          coeffs_126 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_127 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h7f == rs2[7:0]) begin
          coeffs_127 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_128 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h80 == rs2[7:0]) begin
          coeffs_128 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_129 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h81 == rs2[7:0]) begin
          coeffs_129 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_130 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h82 == rs2[7:0]) begin
          coeffs_130 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_131 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h83 == rs2[7:0]) begin
          coeffs_131 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_132 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h84 == rs2[7:0]) begin
          coeffs_132 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_133 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h85 == rs2[7:0]) begin
          coeffs_133 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_134 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h86 == rs2[7:0]) begin
          coeffs_134 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_135 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h87 == rs2[7:0]) begin
          coeffs_135 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_136 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h88 == rs2[7:0]) begin
          coeffs_136 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_137 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h89 == rs2[7:0]) begin
          coeffs_137 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_138 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h8a == rs2[7:0]) begin
          coeffs_138 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_139 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h8b == rs2[7:0]) begin
          coeffs_139 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_140 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h8c == rs2[7:0]) begin
          coeffs_140 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_141 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h8d == rs2[7:0]) begin
          coeffs_141 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_142 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h8e == rs2[7:0]) begin
          coeffs_142 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_143 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h8f == rs2[7:0]) begin
          coeffs_143 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_144 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h90 == rs2[7:0]) begin
          coeffs_144 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_145 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h91 == rs2[7:0]) begin
          coeffs_145 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_146 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h92 == rs2[7:0]) begin
          coeffs_146 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_147 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h93 == rs2[7:0]) begin
          coeffs_147 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_148 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h94 == rs2[7:0]) begin
          coeffs_148 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_149 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h95 == rs2[7:0]) begin
          coeffs_149 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_150 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h96 == rs2[7:0]) begin
          coeffs_150 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_151 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h97 == rs2[7:0]) begin
          coeffs_151 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_152 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h98 == rs2[7:0]) begin
          coeffs_152 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_153 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h99 == rs2[7:0]) begin
          coeffs_153 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_154 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h9a == rs2[7:0]) begin
          coeffs_154 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_155 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h9b == rs2[7:0]) begin
          coeffs_155 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_156 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h9c == rs2[7:0]) begin
          coeffs_156 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_157 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h9d == rs2[7:0]) begin
          coeffs_157 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_158 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h9e == rs2[7:0]) begin
          coeffs_158 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_159 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'h9f == rs2[7:0]) begin
          coeffs_159 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_160 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'ha0 == rs2[7:0]) begin
          coeffs_160 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_161 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'ha1 == rs2[7:0]) begin
          coeffs_161 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_162 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'ha2 == rs2[7:0]) begin
          coeffs_162 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_163 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'ha3 == rs2[7:0]) begin
          coeffs_163 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_164 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'ha4 == rs2[7:0]) begin
          coeffs_164 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_165 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'ha5 == rs2[7:0]) begin
          coeffs_165 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_166 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'ha6 == rs2[7:0]) begin
          coeffs_166 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_167 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'ha7 == rs2[7:0]) begin
          coeffs_167 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_168 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'ha8 == rs2[7:0]) begin
          coeffs_168 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_169 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'ha9 == rs2[7:0]) begin
          coeffs_169 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_170 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'haa == rs2[7:0]) begin
          coeffs_170 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_171 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hab == rs2[7:0]) begin
          coeffs_171 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_172 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hac == rs2[7:0]) begin
          coeffs_172 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_173 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'had == rs2[7:0]) begin
          coeffs_173 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_174 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hae == rs2[7:0]) begin
          coeffs_174 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_175 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'haf == rs2[7:0]) begin
          coeffs_175 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_176 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hb0 == rs2[7:0]) begin
          coeffs_176 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_177 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hb1 == rs2[7:0]) begin
          coeffs_177 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_178 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hb2 == rs2[7:0]) begin
          coeffs_178 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_179 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hb3 == rs2[7:0]) begin
          coeffs_179 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_180 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hb4 == rs2[7:0]) begin
          coeffs_180 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_181 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hb5 == rs2[7:0]) begin
          coeffs_181 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_182 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hb6 == rs2[7:0]) begin
          coeffs_182 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_183 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hb7 == rs2[7:0]) begin
          coeffs_183 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_184 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hb8 == rs2[7:0]) begin
          coeffs_184 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_185 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hb9 == rs2[7:0]) begin
          coeffs_185 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_186 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hba == rs2[7:0]) begin
          coeffs_186 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_187 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hbb == rs2[7:0]) begin
          coeffs_187 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_188 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hbc == rs2[7:0]) begin
          coeffs_188 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_189 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hbd == rs2[7:0]) begin
          coeffs_189 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_190 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hbe == rs2[7:0]) begin
          coeffs_190 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_191 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hbf == rs2[7:0]) begin
          coeffs_191 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_192 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hc0 == rs2[7:0]) begin
          coeffs_192 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_193 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hc1 == rs2[7:0]) begin
          coeffs_193 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_194 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hc2 == rs2[7:0]) begin
          coeffs_194 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_195 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hc3 == rs2[7:0]) begin
          coeffs_195 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_196 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hc4 == rs2[7:0]) begin
          coeffs_196 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_197 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hc5 == rs2[7:0]) begin
          coeffs_197 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_198 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hc6 == rs2[7:0]) begin
          coeffs_198 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_199 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (8'hc7 == rs2[7:0]) begin
          coeffs_199 <= rs1;
        end
      end
    end
    if (reset) begin
      data_0 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_0 <= rs1;
        end
      end
    end
    if (reset) begin
      data_1 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_1 <= data_0;
        end
      end
    end
    if (reset) begin
      data_2 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_2 <= data_1;
        end
      end
    end
    if (reset) begin
      data_3 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_3 <= data_2;
        end
      end
    end
    if (reset) begin
      data_4 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_4 <= data_3;
        end
      end
    end
    if (reset) begin
      data_5 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_5 <= data_4;
        end
      end
    end
    if (reset) begin
      data_6 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_6 <= data_5;
        end
      end
    end
    if (reset) begin
      data_7 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_7 <= data_6;
        end
      end
    end
    if (reset) begin
      data_8 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_8 <= data_7;
        end
      end
    end
    if (reset) begin
      data_9 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_9 <= data_8;
        end
      end
    end
    if (reset) begin
      data_10 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_10 <= data_9;
        end
      end
    end
    if (reset) begin
      data_11 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_11 <= data_10;
        end
      end
    end
    if (reset) begin
      data_12 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_12 <= data_11;
        end
      end
    end
    if (reset) begin
      data_13 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_13 <= data_12;
        end
      end
    end
    if (reset) begin
      data_14 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_14 <= data_13;
        end
      end
    end
    if (reset) begin
      data_15 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_15 <= data_14;
        end
      end
    end
    if (reset) begin
      data_16 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_16 <= data_15;
        end
      end
    end
    if (reset) begin
      data_17 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_17 <= data_16;
        end
      end
    end
    if (reset) begin
      data_18 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_18 <= data_17;
        end
      end
    end
    if (reset) begin
      data_19 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_19 <= data_18;
        end
      end
    end
    if (reset) begin
      data_20 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_20 <= data_19;
        end
      end
    end
    if (reset) begin
      data_21 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_21 <= data_20;
        end
      end
    end
    if (reset) begin
      data_22 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_22 <= data_21;
        end
      end
    end
    if (reset) begin
      data_23 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_23 <= data_22;
        end
      end
    end
    if (reset) begin
      data_24 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_24 <= data_23;
        end
      end
    end
    if (reset) begin
      data_25 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_25 <= data_24;
        end
      end
    end
    if (reset) begin
      data_26 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_26 <= data_25;
        end
      end
    end
    if (reset) begin
      data_27 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_27 <= data_26;
        end
      end
    end
    if (reset) begin
      data_28 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_28 <= data_27;
        end
      end
    end
    if (reset) begin
      data_29 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_29 <= data_28;
        end
      end
    end
    if (reset) begin
      data_30 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_30 <= data_29;
        end
      end
    end
    if (reset) begin
      data_31 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_31 <= data_30;
        end
      end
    end
    if (reset) begin
      data_32 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_32 <= data_31;
        end
      end
    end
    if (reset) begin
      data_33 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_33 <= data_32;
        end
      end
    end
    if (reset) begin
      data_34 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_34 <= data_33;
        end
      end
    end
    if (reset) begin
      data_35 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_35 <= data_34;
        end
      end
    end
    if (reset) begin
      data_36 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_36 <= data_35;
        end
      end
    end
    if (reset) begin
      data_37 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_37 <= data_36;
        end
      end
    end
    if (reset) begin
      data_38 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_38 <= data_37;
        end
      end
    end
    if (reset) begin
      data_39 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_39 <= data_38;
        end
      end
    end
    if (reset) begin
      data_40 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_40 <= data_39;
        end
      end
    end
    if (reset) begin
      data_41 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_41 <= data_40;
        end
      end
    end
    if (reset) begin
      data_42 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_42 <= data_41;
        end
      end
    end
    if (reset) begin
      data_43 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_43 <= data_42;
        end
      end
    end
    if (reset) begin
      data_44 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_44 <= data_43;
        end
      end
    end
    if (reset) begin
      data_45 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_45 <= data_44;
        end
      end
    end
    if (reset) begin
      data_46 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_46 <= data_45;
        end
      end
    end
    if (reset) begin
      data_47 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_47 <= data_46;
        end
      end
    end
    if (reset) begin
      data_48 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_48 <= data_47;
        end
      end
    end
    if (reset) begin
      data_49 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_49 <= data_48;
        end
      end
    end
    if (reset) begin
      data_50 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_50 <= data_49;
        end
      end
    end
    if (reset) begin
      data_51 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_51 <= data_50;
        end
      end
    end
    if (reset) begin
      data_52 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_52 <= data_51;
        end
      end
    end
    if (reset) begin
      data_53 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_53 <= data_52;
        end
      end
    end
    if (reset) begin
      data_54 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_54 <= data_53;
        end
      end
    end
    if (reset) begin
      data_55 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_55 <= data_54;
        end
      end
    end
    if (reset) begin
      data_56 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_56 <= data_55;
        end
      end
    end
    if (reset) begin
      data_57 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_57 <= data_56;
        end
      end
    end
    if (reset) begin
      data_58 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_58 <= data_57;
        end
      end
    end
    if (reset) begin
      data_59 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_59 <= data_58;
        end
      end
    end
    if (reset) begin
      data_60 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_60 <= data_59;
        end
      end
    end
    if (reset) begin
      data_61 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_61 <= data_60;
        end
      end
    end
    if (reset) begin
      data_62 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_62 <= data_61;
        end
      end
    end
    if (reset) begin
      data_63 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_63 <= data_62;
        end
      end
    end
    if (reset) begin
      data_64 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_64 <= data_63;
        end
      end
    end
    if (reset) begin
      data_65 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_65 <= data_64;
        end
      end
    end
    if (reset) begin
      data_66 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_66 <= data_65;
        end
      end
    end
    if (reset) begin
      data_67 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_67 <= data_66;
        end
      end
    end
    if (reset) begin
      data_68 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_68 <= data_67;
        end
      end
    end
    if (reset) begin
      data_69 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_69 <= data_68;
        end
      end
    end
    if (reset) begin
      data_70 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_70 <= data_69;
        end
      end
    end
    if (reset) begin
      data_71 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_71 <= data_70;
        end
      end
    end
    if (reset) begin
      data_72 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_72 <= data_71;
        end
      end
    end
    if (reset) begin
      data_73 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_73 <= data_72;
        end
      end
    end
    if (reset) begin
      data_74 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_74 <= data_73;
        end
      end
    end
    if (reset) begin
      data_75 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_75 <= data_74;
        end
      end
    end
    if (reset) begin
      data_76 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_76 <= data_75;
        end
      end
    end
    if (reset) begin
      data_77 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_77 <= data_76;
        end
      end
    end
    if (reset) begin
      data_78 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_78 <= data_77;
        end
      end
    end
    if (reset) begin
      data_79 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_79 <= data_78;
        end
      end
    end
    if (reset) begin
      data_80 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_80 <= data_79;
        end
      end
    end
    if (reset) begin
      data_81 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_81 <= data_80;
        end
      end
    end
    if (reset) begin
      data_82 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_82 <= data_81;
        end
      end
    end
    if (reset) begin
      data_83 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_83 <= data_82;
        end
      end
    end
    if (reset) begin
      data_84 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_84 <= data_83;
        end
      end
    end
    if (reset) begin
      data_85 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_85 <= data_84;
        end
      end
    end
    if (reset) begin
      data_86 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_86 <= data_85;
        end
      end
    end
    if (reset) begin
      data_87 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_87 <= data_86;
        end
      end
    end
    if (reset) begin
      data_88 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_88 <= data_87;
        end
      end
    end
    if (reset) begin
      data_89 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_89 <= data_88;
        end
      end
    end
    if (reset) begin
      data_90 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_90 <= data_89;
        end
      end
    end
    if (reset) begin
      data_91 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_91 <= data_90;
        end
      end
    end
    if (reset) begin
      data_92 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_92 <= data_91;
        end
      end
    end
    if (reset) begin
      data_93 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_93 <= data_92;
        end
      end
    end
    if (reset) begin
      data_94 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_94 <= data_93;
        end
      end
    end
    if (reset) begin
      data_95 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_95 <= data_94;
        end
      end
    end
    if (reset) begin
      data_96 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_96 <= data_95;
        end
      end
    end
    if (reset) begin
      data_97 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_97 <= data_96;
        end
      end
    end
    if (reset) begin
      data_98 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_98 <= data_97;
        end
      end
    end
    if (reset) begin
      data_99 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_99 <= data_98;
        end
      end
    end
    if (reset) begin
      data_100 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_100 <= data_99;
        end
      end
    end
    if (reset) begin
      data_101 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_101 <= data_100;
        end
      end
    end
    if (reset) begin
      data_102 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_102 <= data_101;
        end
      end
    end
    if (reset) begin
      data_103 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_103 <= data_102;
        end
      end
    end
    if (reset) begin
      data_104 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_104 <= data_103;
        end
      end
    end
    if (reset) begin
      data_105 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_105 <= data_104;
        end
      end
    end
    if (reset) begin
      data_106 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_106 <= data_105;
        end
      end
    end
    if (reset) begin
      data_107 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_107 <= data_106;
        end
      end
    end
    if (reset) begin
      data_108 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_108 <= data_107;
        end
      end
    end
    if (reset) begin
      data_109 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_109 <= data_108;
        end
      end
    end
    if (reset) begin
      data_110 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_110 <= data_109;
        end
      end
    end
    if (reset) begin
      data_111 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_111 <= data_110;
        end
      end
    end
    if (reset) begin
      data_112 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_112 <= data_111;
        end
      end
    end
    if (reset) begin
      data_113 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_113 <= data_112;
        end
      end
    end
    if (reset) begin
      data_114 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_114 <= data_113;
        end
      end
    end
    if (reset) begin
      data_115 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_115 <= data_114;
        end
      end
    end
    if (reset) begin
      data_116 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_116 <= data_115;
        end
      end
    end
    if (reset) begin
      data_117 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_117 <= data_116;
        end
      end
    end
    if (reset) begin
      data_118 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_118 <= data_117;
        end
      end
    end
    if (reset) begin
      data_119 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_119 <= data_118;
        end
      end
    end
    if (reset) begin
      data_120 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_120 <= data_119;
        end
      end
    end
    if (reset) begin
      data_121 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_121 <= data_120;
        end
      end
    end
    if (reset) begin
      data_122 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_122 <= data_121;
        end
      end
    end
    if (reset) begin
      data_123 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_123 <= data_122;
        end
      end
    end
    if (reset) begin
      data_124 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_124 <= data_123;
        end
      end
    end
    if (reset) begin
      data_125 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_125 <= data_124;
        end
      end
    end
    if (reset) begin
      data_126 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_126 <= data_125;
        end
      end
    end
    if (reset) begin
      data_127 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_127 <= data_126;
        end
      end
    end
    if (reset) begin
      data_128 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_128 <= data_127;
        end
      end
    end
    if (reset) begin
      data_129 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_129 <= data_128;
        end
      end
    end
    if (reset) begin
      data_130 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_130 <= data_129;
        end
      end
    end
    if (reset) begin
      data_131 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_131 <= data_130;
        end
      end
    end
    if (reset) begin
      data_132 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_132 <= data_131;
        end
      end
    end
    if (reset) begin
      data_133 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_133 <= data_132;
        end
      end
    end
    if (reset) begin
      data_134 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_134 <= data_133;
        end
      end
    end
    if (reset) begin
      data_135 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_135 <= data_134;
        end
      end
    end
    if (reset) begin
      data_136 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_136 <= data_135;
        end
      end
    end
    if (reset) begin
      data_137 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_137 <= data_136;
        end
      end
    end
    if (reset) begin
      data_138 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_138 <= data_137;
        end
      end
    end
    if (reset) begin
      data_139 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_139 <= data_138;
        end
      end
    end
    if (reset) begin
      data_140 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_140 <= data_139;
        end
      end
    end
    if (reset) begin
      data_141 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_141 <= data_140;
        end
      end
    end
    if (reset) begin
      data_142 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_142 <= data_141;
        end
      end
    end
    if (reset) begin
      data_143 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_143 <= data_142;
        end
      end
    end
    if (reset) begin
      data_144 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_144 <= data_143;
        end
      end
    end
    if (reset) begin
      data_145 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_145 <= data_144;
        end
      end
    end
    if (reset) begin
      data_146 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_146 <= data_145;
        end
      end
    end
    if (reset) begin
      data_147 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_147 <= data_146;
        end
      end
    end
    if (reset) begin
      data_148 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_148 <= data_147;
        end
      end
    end
    if (reset) begin
      data_149 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_149 <= data_148;
        end
      end
    end
    if (reset) begin
      data_150 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_150 <= data_149;
        end
      end
    end
    if (reset) begin
      data_151 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_151 <= data_150;
        end
      end
    end
    if (reset) begin
      data_152 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_152 <= data_151;
        end
      end
    end
    if (reset) begin
      data_153 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_153 <= data_152;
        end
      end
    end
    if (reset) begin
      data_154 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_154 <= data_153;
        end
      end
    end
    if (reset) begin
      data_155 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_155 <= data_154;
        end
      end
    end
    if (reset) begin
      data_156 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_156 <= data_155;
        end
      end
    end
    if (reset) begin
      data_157 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_157 <= data_156;
        end
      end
    end
    if (reset) begin
      data_158 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_158 <= data_157;
        end
      end
    end
    if (reset) begin
      data_159 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_159 <= data_158;
        end
      end
    end
    if (reset) begin
      data_160 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_160 <= data_159;
        end
      end
    end
    if (reset) begin
      data_161 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_161 <= data_160;
        end
      end
    end
    if (reset) begin
      data_162 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_162 <= data_161;
        end
      end
    end
    if (reset) begin
      data_163 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_163 <= data_162;
        end
      end
    end
    if (reset) begin
      data_164 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_164 <= data_163;
        end
      end
    end
    if (reset) begin
      data_165 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_165 <= data_164;
        end
      end
    end
    if (reset) begin
      data_166 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_166 <= data_165;
        end
      end
    end
    if (reset) begin
      data_167 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_167 <= data_166;
        end
      end
    end
    if (reset) begin
      data_168 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_168 <= data_167;
        end
      end
    end
    if (reset) begin
      data_169 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_169 <= data_168;
        end
      end
    end
    if (reset) begin
      data_170 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_170 <= data_169;
        end
      end
    end
    if (reset) begin
      data_171 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_171 <= data_170;
        end
      end
    end
    if (reset) begin
      data_172 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_172 <= data_171;
        end
      end
    end
    if (reset) begin
      data_173 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_173 <= data_172;
        end
      end
    end
    if (reset) begin
      data_174 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_174 <= data_173;
        end
      end
    end
    if (reset) begin
      data_175 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_175 <= data_174;
        end
      end
    end
    if (reset) begin
      data_176 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_176 <= data_175;
        end
      end
    end
    if (reset) begin
      data_177 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_177 <= data_176;
        end
      end
    end
    if (reset) begin
      data_178 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_178 <= data_177;
        end
      end
    end
    if (reset) begin
      data_179 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_179 <= data_178;
        end
      end
    end
    if (reset) begin
      data_180 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_180 <= data_179;
        end
      end
    end
    if (reset) begin
      data_181 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_181 <= data_180;
        end
      end
    end
    if (reset) begin
      data_182 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_182 <= data_181;
        end
      end
    end
    if (reset) begin
      data_183 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_183 <= data_182;
        end
      end
    end
    if (reset) begin
      data_184 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_184 <= data_183;
        end
      end
    end
    if (reset) begin
      data_185 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_185 <= data_184;
        end
      end
    end
    if (reset) begin
      data_186 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_186 <= data_185;
        end
      end
    end
    if (reset) begin
      data_187 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_187 <= data_186;
        end
      end
    end
    if (reset) begin
      data_188 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_188 <= data_187;
        end
      end
    end
    if (reset) begin
      data_189 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_189 <= data_188;
        end
      end
    end
    if (reset) begin
      data_190 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_190 <= data_189;
        end
      end
    end
    if (reset) begin
      data_191 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_191 <= data_190;
        end
      end
    end
    if (reset) begin
      data_192 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_192 <= data_191;
        end
      end
    end
    if (reset) begin
      data_193 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_193 <= data_192;
        end
      end
    end
    if (reset) begin
      data_194 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_194 <= data_193;
        end
      end
    end
    if (reset) begin
      data_195 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_195 <= data_194;
        end
      end
    end
    if (reset) begin
      data_196 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_196 <= data_195;
        end
      end
    end
    if (reset) begin
      data_197 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_197 <= data_196;
        end
      end
    end
    if (reset) begin
      data_198 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_198 <= data_197;
        end
      end
    end
    if (reset) begin
      data_199 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_199 <= data_198;
        end
      end
    end
    if (reset) begin
      result <= 64'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        result <= {{32{_GEN_399[31]}},_GEN_399};
      end else if (insn[6:0] == 7'h2b) begin
        result <= {{32{data_0[31]}},data_0};
      end else begin
        result <= _GEN_400;
      end
    end
  end
endmodule
