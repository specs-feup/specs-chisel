module SCIEPipelined #(parameter XLEN = 32)(
  input         clock,
  input         reset,
  input         valid,
  input  [31:0] insn,
  input  [31:0] rs1,
  input  [31:0] rs2,
  output [31:0] rd
);
  reg [31:0] coeffs_0;
  reg [31:0] coeffs_1;
  reg [31:0] coeffs_2;
  reg [31:0] coeffs_3;
  reg [31:0] coeffs_4;
  reg [31:0] coeffs_5;
  reg [31:0] coeffs_6;
  reg [31:0] coeffs_7;
  reg [31:0] coeffs_8;
  reg [31:0] coeffs_9;
  reg [31:0] coeffs_10;
  reg [31:0] coeffs_11;
  reg [31:0] coeffs_12;
  reg [31:0] coeffs_13;
  reg [31:0] coeffs_14;
  reg [31:0] coeffs_15;
  reg [31:0] coeffs_16;
  reg [31:0] coeffs_17;
  reg [31:0] coeffs_18;
  reg [31:0] coeffs_19;
  reg [31:0] coeffs_20;
  reg [31:0] coeffs_21;
  reg [31:0] coeffs_22;
  reg [31:0] coeffs_23;
  reg [31:0] coeffs_24;
  reg [31:0] coeffs_25;
  reg [31:0] coeffs_26;
  reg [31:0] coeffs_27;
  reg [31:0] coeffs_28;
  reg [31:0] coeffs_29;
  reg [31:0] coeffs_30;
  reg [31:0] coeffs_31;
  reg [31:0] coeffs_32;
  reg [31:0] coeffs_33;
  reg [31:0] coeffs_34;
  reg [31:0] coeffs_35;
  reg [31:0] coeffs_36;
  reg [31:0] coeffs_37;
  reg [31:0] coeffs_38;
  reg [31:0] coeffs_39;
  reg [31:0] coeffs_40;
  reg [31:0] coeffs_41;
  reg [31:0] coeffs_42;
  reg [31:0] coeffs_43;
  reg [31:0] coeffs_44;
  reg [31:0] coeffs_45;
  reg [31:0] coeffs_46;
  reg [31:0] coeffs_47;
  reg [31:0] coeffs_48;
  reg [31:0] coeffs_49;
  reg [31:0] coeffs_50;
  reg [31:0] coeffs_51;
  reg [31:0] coeffs_52;
  reg [31:0] coeffs_53;
  reg [31:0] coeffs_54;
  reg [31:0] coeffs_55;
  reg [31:0] coeffs_56;
  reg [31:0] coeffs_57;
  reg [31:0] coeffs_58;
  reg [31:0] coeffs_59;
  reg [31:0] coeffs_60;
  reg [31:0] coeffs_61;
  reg [31:0] coeffs_62;
  reg [31:0] coeffs_63;
  reg [31:0] coeffs_64;
  reg [31:0] coeffs_65;
  reg [31:0] coeffs_66;
  reg [31:0] coeffs_67;
  reg [31:0] coeffs_68;
  reg [31:0] coeffs_69;
  reg [31:0] coeffs_70;
  reg [31:0] coeffs_71;
  reg [31:0] coeffs_72;
  reg [31:0] coeffs_73;
  reg [31:0] coeffs_74;
  reg [31:0] coeffs_75;
  reg [31:0] coeffs_76;
  reg [31:0] coeffs_77;
  reg [31:0] coeffs_78;
  reg [31:0] coeffs_79;
  reg [31:0] coeffs_80;
  reg [31:0] coeffs_81;
  reg [31:0] coeffs_82;
  reg [31:0] coeffs_83;
  reg [31:0] coeffs_84;
  reg [31:0] coeffs_85;
  reg [31:0] coeffs_86;
  reg [31:0] coeffs_87;
  reg [31:0] coeffs_88;
  reg [31:0] coeffs_89;
  reg [31:0] coeffs_90;
  reg [31:0] coeffs_91;
  reg [31:0] coeffs_92;
  reg [31:0] coeffs_93;
  reg [31:0] coeffs_94;
  reg [31:0] coeffs_95;
  reg [31:0] coeffs_96;
  reg [31:0] coeffs_97;
  reg [31:0] coeffs_98;
  reg [31:0] coeffs_99;
  reg [31:0] coeffs_100;
  reg [31:0] coeffs_101;
  reg [31:0] coeffs_102;
  reg [31:0] coeffs_103;
  reg [31:0] coeffs_104;
  reg [31:0] coeffs_105;
  reg [31:0] coeffs_106;
  reg [31:0] coeffs_107;
  reg [31:0] coeffs_108;
  reg [31:0] coeffs_109;
  reg [31:0] coeffs_110;
  reg [31:0] coeffs_111;
  reg [31:0] coeffs_112;
  reg [31:0] coeffs_113;
  reg [31:0] coeffs_114;
  reg [31:0] coeffs_115;
  reg [31:0] coeffs_116;
  reg [31:0] coeffs_117;
  reg [31:0] coeffs_118;
  reg [31:0] coeffs_119;
  reg [31:0] coeffs_120;
  reg [31:0] coeffs_121;
  reg [31:0] coeffs_122;
  reg [31:0] coeffs_123;
  reg [31:0] coeffs_124;
  reg [31:0] coeffs_125;
  reg [31:0] coeffs_126;
  reg [31:0] coeffs_127;
  reg [31:0] coeffs_128;
  reg [31:0] coeffs_129;
  reg [31:0] coeffs_130;
  reg [31:0] coeffs_131;
  reg [31:0] coeffs_132;
  reg [31:0] coeffs_133;
  reg [31:0] coeffs_134;
  reg [31:0] coeffs_135;
  reg [31:0] coeffs_136;
  reg [31:0] coeffs_137;
  reg [31:0] coeffs_138;
  reg [31:0] coeffs_139;
  reg [31:0] coeffs_140;
  reg [31:0] coeffs_141;
  reg [31:0] coeffs_142;
  reg [31:0] coeffs_143;
  reg [31:0] coeffs_144;
  reg [31:0] coeffs_145;
  reg [31:0] coeffs_146;
  reg [31:0] coeffs_147;
  reg [31:0] coeffs_148;
  reg [31:0] coeffs_149;
  reg [31:0] coeffs_150;
  reg [31:0] coeffs_151;
  reg [31:0] coeffs_152;
  reg [31:0] coeffs_153;
  reg [31:0] coeffs_154;
  reg [31:0] coeffs_155;
  reg [31:0] coeffs_156;
  reg [31:0] coeffs_157;
  reg [31:0] coeffs_158;
  reg [31:0] coeffs_159;
  reg [31:0] coeffs_160;
  reg [31:0] coeffs_161;
  reg [31:0] coeffs_162;
  reg [31:0] coeffs_163;
  reg [31:0] coeffs_164;
  reg [31:0] coeffs_165;
  reg [31:0] coeffs_166;
  reg [31:0] coeffs_167;
  reg [31:0] coeffs_168;
  reg [31:0] coeffs_169;
  reg [31:0] coeffs_170;
  reg [31:0] coeffs_171;
  reg [31:0] coeffs_172;
  reg [31:0] coeffs_173;
  reg [31:0] coeffs_174;
  reg [31:0] coeffs_175;
  reg [31:0] coeffs_176;
  reg [31:0] coeffs_177;
  reg [31:0] coeffs_178;
  reg [31:0] coeffs_179;
  reg [31:0] coeffs_180;
  reg [31:0] coeffs_181;
  reg [31:0] coeffs_182;
  reg [31:0] coeffs_183;
  reg [31:0] coeffs_184;
  reg [31:0] coeffs_185;
  reg [31:0] coeffs_186;
  reg [31:0] coeffs_187;
  reg [31:0] coeffs_188;
  reg [31:0] coeffs_189;
  reg [31:0] coeffs_190;
  reg [31:0] coeffs_191;
  reg [31:0] coeffs_192;
  reg [31:0] coeffs_193;
  reg [31:0] coeffs_194;
  reg [31:0] coeffs_195;
  reg [31:0] coeffs_196;
  reg [31:0] coeffs_197;
  reg [31:0] coeffs_198;
  reg [31:0] coeffs_199;
  reg [31:0] coeffs_200;
  reg [31:0] coeffs_201;
  reg [31:0] coeffs_202;
  reg [31:0] coeffs_203;
  reg [31:0] coeffs_204;
  reg [31:0] coeffs_205;
  reg [31:0] coeffs_206;
  reg [31:0] coeffs_207;
  reg [31:0] coeffs_208;
  reg [31:0] coeffs_209;
  reg [31:0] coeffs_210;
  reg [31:0] coeffs_211;
  reg [31:0] coeffs_212;
  reg [31:0] coeffs_213;
  reg [31:0] coeffs_214;
  reg [31:0] coeffs_215;
  reg [31:0] coeffs_216;
  reg [31:0] coeffs_217;
  reg [31:0] coeffs_218;
  reg [31:0] coeffs_219;
  reg [31:0] coeffs_220;
  reg [31:0] coeffs_221;
  reg [31:0] coeffs_222;
  reg [31:0] coeffs_223;
  reg [31:0] coeffs_224;
  reg [31:0] coeffs_225;
  reg [31:0] coeffs_226;
  reg [31:0] coeffs_227;
  reg [31:0] coeffs_228;
  reg [31:0] coeffs_229;
  reg [31:0] coeffs_230;
  reg [31:0] coeffs_231;
  reg [31:0] coeffs_232;
  reg [31:0] coeffs_233;
  reg [31:0] coeffs_234;
  reg [31:0] coeffs_235;
  reg [31:0] coeffs_236;
  reg [31:0] coeffs_237;
  reg [31:0] coeffs_238;
  reg [31:0] coeffs_239;
  reg [31:0] coeffs_240;
  reg [31:0] coeffs_241;
  reg [31:0] coeffs_242;
  reg [31:0] coeffs_243;
  reg [31:0] coeffs_244;
  reg [31:0] coeffs_245;
  reg [31:0] coeffs_246;
  reg [31:0] coeffs_247;
  reg [31:0] coeffs_248;
  reg [31:0] coeffs_249;
  reg [31:0] coeffs_250;
  reg [31:0] coeffs_251;
  reg [31:0] coeffs_252;
  reg [31:0] coeffs_253;
  reg [31:0] coeffs_254;
  reg [31:0] coeffs_255;
  reg [31:0] coeffs_256;
  reg [31:0] coeffs_257;
  reg [31:0] coeffs_258;
  reg [31:0] coeffs_259;
  reg [31:0] coeffs_260;
  reg [31:0] coeffs_261;
  reg [31:0] coeffs_262;
  reg [31:0] coeffs_263;
  reg [31:0] coeffs_264;
  reg [31:0] coeffs_265;
  reg [31:0] coeffs_266;
  reg [31:0] coeffs_267;
  reg [31:0] coeffs_268;
  reg [31:0] coeffs_269;
  reg [31:0] coeffs_270;
  reg [31:0] coeffs_271;
  reg [31:0] coeffs_272;
  reg [31:0] coeffs_273;
  reg [31:0] coeffs_274;
  reg [31:0] coeffs_275;
  reg [31:0] coeffs_276;
  reg [31:0] coeffs_277;
  reg [31:0] coeffs_278;
  reg [31:0] coeffs_279;
  reg [31:0] coeffs_280;
  reg [31:0] coeffs_281;
  reg [31:0] coeffs_282;
  reg [31:0] coeffs_283;
  reg [31:0] coeffs_284;
  reg [31:0] coeffs_285;
  reg [31:0] coeffs_286;
  reg [31:0] coeffs_287;
  reg [31:0] coeffs_288;
  reg [31:0] coeffs_289;
  reg [31:0] coeffs_290;
  reg [31:0] coeffs_291;
  reg [31:0] coeffs_292;
  reg [31:0] coeffs_293;
  reg [31:0] coeffs_294;
  reg [31:0] coeffs_295;
  reg [31:0] coeffs_296;
  reg [31:0] coeffs_297;
  reg [31:0] coeffs_298;
  reg [31:0] coeffs_299;
  reg [31:0] coeffs_300;
  reg [31:0] coeffs_301;
  reg [31:0] coeffs_302;
  reg [31:0] coeffs_303;
  reg [31:0] coeffs_304;
  reg [31:0] coeffs_305;
  reg [31:0] coeffs_306;
  reg [31:0] coeffs_307;
  reg [31:0] coeffs_308;
  reg [31:0] coeffs_309;
  reg [31:0] coeffs_310;
  reg [31:0] coeffs_311;
  reg [31:0] coeffs_312;
  reg [31:0] coeffs_313;
  reg [31:0] coeffs_314;
  reg [31:0] coeffs_315;
  reg [31:0] coeffs_316;
  reg [31:0] coeffs_317;
  reg [31:0] coeffs_318;
  reg [31:0] coeffs_319;
  reg [31:0] coeffs_320;
  reg [31:0] coeffs_321;
  reg [31:0] coeffs_322;
  reg [31:0] coeffs_323;
  reg [31:0] coeffs_324;
  reg [31:0] coeffs_325;
  reg [31:0] coeffs_326;
  reg [31:0] coeffs_327;
  reg [31:0] coeffs_328;
  reg [31:0] coeffs_329;
  reg [31:0] coeffs_330;
  reg [31:0] coeffs_331;
  reg [31:0] coeffs_332;
  reg [31:0] coeffs_333;
  reg [31:0] coeffs_334;
  reg [31:0] coeffs_335;
  reg [31:0] coeffs_336;
  reg [31:0] coeffs_337;
  reg [31:0] coeffs_338;
  reg [31:0] coeffs_339;
  reg [31:0] coeffs_340;
  reg [31:0] coeffs_341;
  reg [31:0] coeffs_342;
  reg [31:0] coeffs_343;
  reg [31:0] coeffs_344;
  reg [31:0] coeffs_345;
  reg [31:0] coeffs_346;
  reg [31:0] coeffs_347;
  reg [31:0] coeffs_348;
  reg [31:0] coeffs_349;
  reg [31:0] coeffs_350;
  reg [31:0] coeffs_351;
  reg [31:0] coeffs_352;
  reg [31:0] coeffs_353;
  reg [31:0] coeffs_354;
  reg [31:0] coeffs_355;
  reg [31:0] coeffs_356;
  reg [31:0] coeffs_357;
  reg [31:0] coeffs_358;
  reg [31:0] coeffs_359;
  reg [31:0] coeffs_360;
  reg [31:0] coeffs_361;
  reg [31:0] coeffs_362;
  reg [31:0] coeffs_363;
  reg [31:0] coeffs_364;
  reg [31:0] coeffs_365;
  reg [31:0] coeffs_366;
  reg [31:0] coeffs_367;
  reg [31:0] coeffs_368;
  reg [31:0] coeffs_369;
  reg [31:0] coeffs_370;
  reg [31:0] coeffs_371;
  reg [31:0] coeffs_372;
  reg [31:0] coeffs_373;
  reg [31:0] coeffs_374;
  reg [31:0] coeffs_375;
  reg [31:0] coeffs_376;
  reg [31:0] coeffs_377;
  reg [31:0] coeffs_378;
  reg [31:0] coeffs_379;
  reg [31:0] coeffs_380;
  reg [31:0] coeffs_381;
  reg [31:0] coeffs_382;
  reg [31:0] coeffs_383;
  reg [31:0] coeffs_384;
  reg [31:0] coeffs_385;
  reg [31:0] coeffs_386;
  reg [31:0] coeffs_387;
  reg [31:0] coeffs_388;
  reg [31:0] coeffs_389;
  reg [31:0] coeffs_390;
  reg [31:0] coeffs_391;
  reg [31:0] coeffs_392;
  reg [31:0] coeffs_393;
  reg [31:0] coeffs_394;
  reg [31:0] coeffs_395;
  reg [31:0] coeffs_396;
  reg [31:0] coeffs_397;
  reg [31:0] coeffs_398;
  reg [31:0] coeffs_399;
  reg [31:0] coeffs_400;
  reg [31:0] coeffs_401;
  reg [31:0] coeffs_402;
  reg [31:0] coeffs_403;
  reg [31:0] coeffs_404;
  reg [31:0] coeffs_405;
  reg [31:0] coeffs_406;
  reg [31:0] coeffs_407;
  reg [31:0] coeffs_408;
  reg [31:0] coeffs_409;
  reg [31:0] coeffs_410;
  reg [31:0] coeffs_411;
  reg [31:0] coeffs_412;
  reg [31:0] coeffs_413;
  reg [31:0] coeffs_414;
  reg [31:0] coeffs_415;
  reg [31:0] coeffs_416;
  reg [31:0] coeffs_417;
  reg [31:0] coeffs_418;
  reg [31:0] coeffs_419;
  reg [31:0] coeffs_420;
  reg [31:0] coeffs_421;
  reg [31:0] coeffs_422;
  reg [31:0] coeffs_423;
  reg [31:0] coeffs_424;
  reg [31:0] coeffs_425;
  reg [31:0] coeffs_426;
  reg [31:0] coeffs_427;
  reg [31:0] coeffs_428;
  reg [31:0] coeffs_429;
  reg [31:0] coeffs_430;
  reg [31:0] coeffs_431;
  reg [31:0] coeffs_432;
  reg [31:0] coeffs_433;
  reg [31:0] coeffs_434;
  reg [31:0] coeffs_435;
  reg [31:0] coeffs_436;
  reg [31:0] coeffs_437;
  reg [31:0] coeffs_438;
  reg [31:0] coeffs_439;
  reg [31:0] coeffs_440;
  reg [31:0] coeffs_441;
  reg [31:0] coeffs_442;
  reg [31:0] coeffs_443;
  reg [31:0] coeffs_444;
  reg [31:0] coeffs_445;
  reg [31:0] coeffs_446;
  reg [31:0] coeffs_447;
  reg [31:0] coeffs_448;
  reg [31:0] coeffs_449;
  reg [31:0] coeffs_450;
  reg [31:0] coeffs_451;
  reg [31:0] coeffs_452;
  reg [31:0] coeffs_453;
  reg [31:0] coeffs_454;
  reg [31:0] coeffs_455;
  reg [31:0] coeffs_456;
  reg [31:0] coeffs_457;
  reg [31:0] coeffs_458;
  reg [31:0] coeffs_459;
  reg [31:0] coeffs_460;
  reg [31:0] coeffs_461;
  reg [31:0] coeffs_462;
  reg [31:0] coeffs_463;
  reg [31:0] coeffs_464;
  reg [31:0] coeffs_465;
  reg [31:0] coeffs_466;
  reg [31:0] coeffs_467;
  reg [31:0] coeffs_468;
  reg [31:0] coeffs_469;
  reg [31:0] coeffs_470;
  reg [31:0] coeffs_471;
  reg [31:0] coeffs_472;
  reg [31:0] coeffs_473;
  reg [31:0] coeffs_474;
  reg [31:0] coeffs_475;
  reg [31:0] coeffs_476;
  reg [31:0] coeffs_477;
  reg [31:0] coeffs_478;
  reg [31:0] coeffs_479;
  reg [31:0] coeffs_480;
  reg [31:0] coeffs_481;
  reg [31:0] coeffs_482;
  reg [31:0] coeffs_483;
  reg [31:0] coeffs_484;
  reg [31:0] coeffs_485;
  reg [31:0] coeffs_486;
  reg [31:0] coeffs_487;
  reg [31:0] coeffs_488;
  reg [31:0] coeffs_489;
  reg [31:0] coeffs_490;
  reg [31:0] coeffs_491;
  reg [31:0] coeffs_492;
  reg [31:0] coeffs_493;
  reg [31:0] coeffs_494;
  reg [31:0] coeffs_495;
  reg [31:0] coeffs_496;
  reg [31:0] coeffs_497;
  reg [31:0] coeffs_498;
  reg [31:0] coeffs_499;
  reg [31:0] data_0;
  reg [31:0] data_1;
  reg [31:0] data_2;
  reg [31:0] data_3;
  reg [31:0] data_4;
  reg [31:0] data_5;
  reg [31:0] data_6;
  reg [31:0] data_7;
  reg [31:0] data_8;
  reg [31:0] data_9;
  reg [31:0] data_10;
  reg [31:0] data_11;
  reg [31:0] data_12;
  reg [31:0] data_13;
  reg [31:0] data_14;
  reg [31:0] data_15;
  reg [31:0] data_16;
  reg [31:0] data_17;
  reg [31:0] data_18;
  reg [31:0] data_19;
  reg [31:0] data_20;
  reg [31:0] data_21;
  reg [31:0] data_22;
  reg [31:0] data_23;
  reg [31:0] data_24;
  reg [31:0] data_25;
  reg [31:0] data_26;
  reg [31:0] data_27;
  reg [31:0] data_28;
  reg [31:0] data_29;
  reg [31:0] data_30;
  reg [31:0] data_31;
  reg [31:0] data_32;
  reg [31:0] data_33;
  reg [31:0] data_34;
  reg [31:0] data_35;
  reg [31:0] data_36;
  reg [31:0] data_37;
  reg [31:0] data_38;
  reg [31:0] data_39;
  reg [31:0] data_40;
  reg [31:0] data_41;
  reg [31:0] data_42;
  reg [31:0] data_43;
  reg [31:0] data_44;
  reg [31:0] data_45;
  reg [31:0] data_46;
  reg [31:0] data_47;
  reg [31:0] data_48;
  reg [31:0] data_49;
  reg [31:0] data_50;
  reg [31:0] data_51;
  reg [31:0] data_52;
  reg [31:0] data_53;
  reg [31:0] data_54;
  reg [31:0] data_55;
  reg [31:0] data_56;
  reg [31:0] data_57;
  reg [31:0] data_58;
  reg [31:0] data_59;
  reg [31:0] data_60;
  reg [31:0] data_61;
  reg [31:0] data_62;
  reg [31:0] data_63;
  reg [31:0] data_64;
  reg [31:0] data_65;
  reg [31:0] data_66;
  reg [31:0] data_67;
  reg [31:0] data_68;
  reg [31:0] data_69;
  reg [31:0] data_70;
  reg [31:0] data_71;
  reg [31:0] data_72;
  reg [31:0] data_73;
  reg [31:0] data_74;
  reg [31:0] data_75;
  reg [31:0] data_76;
  reg [31:0] data_77;
  reg [31:0] data_78;
  reg [31:0] data_79;
  reg [31:0] data_80;
  reg [31:0] data_81;
  reg [31:0] data_82;
  reg [31:0] data_83;
  reg [31:0] data_84;
  reg [31:0] data_85;
  reg [31:0] data_86;
  reg [31:0] data_87;
  reg [31:0] data_88;
  reg [31:0] data_89;
  reg [31:0] data_90;
  reg [31:0] data_91;
  reg [31:0] data_92;
  reg [31:0] data_93;
  reg [31:0] data_94;
  reg [31:0] data_95;
  reg [31:0] data_96;
  reg [31:0] data_97;
  reg [31:0] data_98;
  reg [31:0] data_99;
  reg [31:0] data_100;
  reg [31:0] data_101;
  reg [31:0] data_102;
  reg [31:0] data_103;
  reg [31:0] data_104;
  reg [31:0] data_105;
  reg [31:0] data_106;
  reg [31:0] data_107;
  reg [31:0] data_108;
  reg [31:0] data_109;
  reg [31:0] data_110;
  reg [31:0] data_111;
  reg [31:0] data_112;
  reg [31:0] data_113;
  reg [31:0] data_114;
  reg [31:0] data_115;
  reg [31:0] data_116;
  reg [31:0] data_117;
  reg [31:0] data_118;
  reg [31:0] data_119;
  reg [31:0] data_120;
  reg [31:0] data_121;
  reg [31:0] data_122;
  reg [31:0] data_123;
  reg [31:0] data_124;
  reg [31:0] data_125;
  reg [31:0] data_126;
  reg [31:0] data_127;
  reg [31:0] data_128;
  reg [31:0] data_129;
  reg [31:0] data_130;
  reg [31:0] data_131;
  reg [31:0] data_132;
  reg [31:0] data_133;
  reg [31:0] data_134;
  reg [31:0] data_135;
  reg [31:0] data_136;
  reg [31:0] data_137;
  reg [31:0] data_138;
  reg [31:0] data_139;
  reg [31:0] data_140;
  reg [31:0] data_141;
  reg [31:0] data_142;
  reg [31:0] data_143;
  reg [31:0] data_144;
  reg [31:0] data_145;
  reg [31:0] data_146;
  reg [31:0] data_147;
  reg [31:0] data_148;
  reg [31:0] data_149;
  reg [31:0] data_150;
  reg [31:0] data_151;
  reg [31:0] data_152;
  reg [31:0] data_153;
  reg [31:0] data_154;
  reg [31:0] data_155;
  reg [31:0] data_156;
  reg [31:0] data_157;
  reg [31:0] data_158;
  reg [31:0] data_159;
  reg [31:0] data_160;
  reg [31:0] data_161;
  reg [31:0] data_162;
  reg [31:0] data_163;
  reg [31:0] data_164;
  reg [31:0] data_165;
  reg [31:0] data_166;
  reg [31:0] data_167;
  reg [31:0] data_168;
  reg [31:0] data_169;
  reg [31:0] data_170;
  reg [31:0] data_171;
  reg [31:0] data_172;
  reg [31:0] data_173;
  reg [31:0] data_174;
  reg [31:0] data_175;
  reg [31:0] data_176;
  reg [31:0] data_177;
  reg [31:0] data_178;
  reg [31:0] data_179;
  reg [31:0] data_180;
  reg [31:0] data_181;
  reg [31:0] data_182;
  reg [31:0] data_183;
  reg [31:0] data_184;
  reg [31:0] data_185;
  reg [31:0] data_186;
  reg [31:0] data_187;
  reg [31:0] data_188;
  reg [31:0] data_189;
  reg [31:0] data_190;
  reg [31:0] data_191;
  reg [31:0] data_192;
  reg [31:0] data_193;
  reg [31:0] data_194;
  reg [31:0] data_195;
  reg [31:0] data_196;
  reg [31:0] data_197;
  reg [31:0] data_198;
  reg [31:0] data_199;
  reg [31:0] data_200;
  reg [31:0] data_201;
  reg [31:0] data_202;
  reg [31:0] data_203;
  reg [31:0] data_204;
  reg [31:0] data_205;
  reg [31:0] data_206;
  reg [31:0] data_207;
  reg [31:0] data_208;
  reg [31:0] data_209;
  reg [31:0] data_210;
  reg [31:0] data_211;
  reg [31:0] data_212;
  reg [31:0] data_213;
  reg [31:0] data_214;
  reg [31:0] data_215;
  reg [31:0] data_216;
  reg [31:0] data_217;
  reg [31:0] data_218;
  reg [31:0] data_219;
  reg [31:0] data_220;
  reg [31:0] data_221;
  reg [31:0] data_222;
  reg [31:0] data_223;
  reg [31:0] data_224;
  reg [31:0] data_225;
  reg [31:0] data_226;
  reg [31:0] data_227;
  reg [31:0] data_228;
  reg [31:0] data_229;
  reg [31:0] data_230;
  reg [31:0] data_231;
  reg [31:0] data_232;
  reg [31:0] data_233;
  reg [31:0] data_234;
  reg [31:0] data_235;
  reg [31:0] data_236;
  reg [31:0] data_237;
  reg [31:0] data_238;
  reg [31:0] data_239;
  reg [31:0] data_240;
  reg [31:0] data_241;
  reg [31:0] data_242;
  reg [31:0] data_243;
  reg [31:0] data_244;
  reg [31:0] data_245;
  reg [31:0] data_246;
  reg [31:0] data_247;
  reg [31:0] data_248;
  reg [31:0] data_249;
  reg [31:0] data_250;
  reg [31:0] data_251;
  reg [31:0] data_252;
  reg [31:0] data_253;
  reg [31:0] data_254;
  reg [31:0] data_255;
  reg [31:0] data_256;
  reg [31:0] data_257;
  reg [31:0] data_258;
  reg [31:0] data_259;
  reg [31:0] data_260;
  reg [31:0] data_261;
  reg [31:0] data_262;
  reg [31:0] data_263;
  reg [31:0] data_264;
  reg [31:0] data_265;
  reg [31:0] data_266;
  reg [31:0] data_267;
  reg [31:0] data_268;
  reg [31:0] data_269;
  reg [31:0] data_270;
  reg [31:0] data_271;
  reg [31:0] data_272;
  reg [31:0] data_273;
  reg [31:0] data_274;
  reg [31:0] data_275;
  reg [31:0] data_276;
  reg [31:0] data_277;
  reg [31:0] data_278;
  reg [31:0] data_279;
  reg [31:0] data_280;
  reg [31:0] data_281;
  reg [31:0] data_282;
  reg [31:0] data_283;
  reg [31:0] data_284;
  reg [31:0] data_285;
  reg [31:0] data_286;
  reg [31:0] data_287;
  reg [31:0] data_288;
  reg [31:0] data_289;
  reg [31:0] data_290;
  reg [31:0] data_291;
  reg [31:0] data_292;
  reg [31:0] data_293;
  reg [31:0] data_294;
  reg [31:0] data_295;
  reg [31:0] data_296;
  reg [31:0] data_297;
  reg [31:0] data_298;
  reg [31:0] data_299;
  reg [31:0] data_300;
  reg [31:0] data_301;
  reg [31:0] data_302;
  reg [31:0] data_303;
  reg [31:0] data_304;
  reg [31:0] data_305;
  reg [31:0] data_306;
  reg [31:0] data_307;
  reg [31:0] data_308;
  reg [31:0] data_309;
  reg [31:0] data_310;
  reg [31:0] data_311;
  reg [31:0] data_312;
  reg [31:0] data_313;
  reg [31:0] data_314;
  reg [31:0] data_315;
  reg [31:0] data_316;
  reg [31:0] data_317;
  reg [31:0] data_318;
  reg [31:0] data_319;
  reg [31:0] data_320;
  reg [31:0] data_321;
  reg [31:0] data_322;
  reg [31:0] data_323;
  reg [31:0] data_324;
  reg [31:0] data_325;
  reg [31:0] data_326;
  reg [31:0] data_327;
  reg [31:0] data_328;
  reg [31:0] data_329;
  reg [31:0] data_330;
  reg [31:0] data_331;
  reg [31:0] data_332;
  reg [31:0] data_333;
  reg [31:0] data_334;
  reg [31:0] data_335;
  reg [31:0] data_336;
  reg [31:0] data_337;
  reg [31:0] data_338;
  reg [31:0] data_339;
  reg [31:0] data_340;
  reg [31:0] data_341;
  reg [31:0] data_342;
  reg [31:0] data_343;
  reg [31:0] data_344;
  reg [31:0] data_345;
  reg [31:0] data_346;
  reg [31:0] data_347;
  reg [31:0] data_348;
  reg [31:0] data_349;
  reg [31:0] data_350;
  reg [31:0] data_351;
  reg [31:0] data_352;
  reg [31:0] data_353;
  reg [31:0] data_354;
  reg [31:0] data_355;
  reg [31:0] data_356;
  reg [31:0] data_357;
  reg [31:0] data_358;
  reg [31:0] data_359;
  reg [31:0] data_360;
  reg [31:0] data_361;
  reg [31:0] data_362;
  reg [31:0] data_363;
  reg [31:0] data_364;
  reg [31:0] data_365;
  reg [31:0] data_366;
  reg [31:0] data_367;
  reg [31:0] data_368;
  reg [31:0] data_369;
  reg [31:0] data_370;
  reg [31:0] data_371;
  reg [31:0] data_372;
  reg [31:0] data_373;
  reg [31:0] data_374;
  reg [31:0] data_375;
  reg [31:0] data_376;
  reg [31:0] data_377;
  reg [31:0] data_378;
  reg [31:0] data_379;
  reg [31:0] data_380;
  reg [31:0] data_381;
  reg [31:0] data_382;
  reg [31:0] data_383;
  reg [31:0] data_384;
  reg [31:0] data_385;
  reg [31:0] data_386;
  reg [31:0] data_387;
  reg [31:0] data_388;
  reg [31:0] data_389;
  reg [31:0] data_390;
  reg [31:0] data_391;
  reg [31:0] data_392;
  reg [31:0] data_393;
  reg [31:0] data_394;
  reg [31:0] data_395;
  reg [31:0] data_396;
  reg [31:0] data_397;
  reg [31:0] data_398;
  reg [31:0] data_399;
  reg [31:0] data_400;
  reg [31:0] data_401;
  reg [31:0] data_402;
  reg [31:0] data_403;
  reg [31:0] data_404;
  reg [31:0] data_405;
  reg [31:0] data_406;
  reg [31:0] data_407;
  reg [31:0] data_408;
  reg [31:0] data_409;
  reg [31:0] data_410;
  reg [31:0] data_411;
  reg [31:0] data_412;
  reg [31:0] data_413;
  reg [31:0] data_414;
  reg [31:0] data_415;
  reg [31:0] data_416;
  reg [31:0] data_417;
  reg [31:0] data_418;
  reg [31:0] data_419;
  reg [31:0] data_420;
  reg [31:0] data_421;
  reg [31:0] data_422;
  reg [31:0] data_423;
  reg [31:0] data_424;
  reg [31:0] data_425;
  reg [31:0] data_426;
  reg [31:0] data_427;
  reg [31:0] data_428;
  reg [31:0] data_429;
  reg [31:0] data_430;
  reg [31:0] data_431;
  reg [31:0] data_432;
  reg [31:0] data_433;
  reg [31:0] data_434;
  reg [31:0] data_435;
  reg [31:0] data_436;
  reg [31:0] data_437;
  reg [31:0] data_438;
  reg [31:0] data_439;
  reg [31:0] data_440;
  reg [31:0] data_441;
  reg [31:0] data_442;
  reg [31:0] data_443;
  reg [31:0] data_444;
  reg [31:0] data_445;
  reg [31:0] data_446;
  reg [31:0] data_447;
  reg [31:0] data_448;
  reg [31:0] data_449;
  reg [31:0] data_450;
  reg [31:0] data_451;
  reg [31:0] data_452;
  reg [31:0] data_453;
  reg [31:0] data_454;
  reg [31:0] data_455;
  reg [31:0] data_456;
  reg [31:0] data_457;
  reg [31:0] data_458;
  reg [31:0] data_459;
  reg [31:0] data_460;
  reg [31:0] data_461;
  reg [31:0] data_462;
  reg [31:0] data_463;
  reg [31:0] data_464;
  reg [31:0] data_465;
  reg [31:0] data_466;
  reg [31:0] data_467;
  reg [31:0] data_468;
  reg [31:0] data_469;
  reg [31:0] data_470;
  reg [31:0] data_471;
  reg [31:0] data_472;
  reg [31:0] data_473;
  reg [31:0] data_474;
  reg [31:0] data_475;
  reg [31:0] data_476;
  reg [31:0] data_477;
  reg [31:0] data_478;
  reg [31:0] data_479;
  reg [31:0] data_480;
  reg [31:0] data_481;
  reg [31:0] data_482;
  reg [31:0] data_483;
  reg [31:0] data_484;
  reg [31:0] data_485;
  reg [31:0] data_486;
  reg [31:0] data_487;
  reg [31:0] data_488;
  reg [31:0] data_489;
  reg [31:0] data_490;
  reg [31:0] data_491;
  reg [31:0] data_492;
  reg [31:0] data_493;
  reg [31:0] data_494;
  reg [31:0] data_495;
  reg [31:0] data_496;
  reg [31:0] data_497;
  reg [31:0] data_498;
  reg [31:0] data_499;
  reg [63:0] result;
  wire [31:0] _GEN_501 = 9'h1 == rs2[8:0] ? coeffs_1 : coeffs_0;
  wire [31:0] _GEN_502 = 9'h2 == rs2[8:0] ? coeffs_2 : _GEN_501;
  wire [31:0] _GEN_503 = 9'h3 == rs2[8:0] ? coeffs_3 : _GEN_502;
  wire [31:0] _GEN_504 = 9'h4 == rs2[8:0] ? coeffs_4 : _GEN_503;
  wire [31:0] _GEN_505 = 9'h5 == rs2[8:0] ? coeffs_5 : _GEN_504;
  wire [31:0] _GEN_506 = 9'h6 == rs2[8:0] ? coeffs_6 : _GEN_505;
  wire [31:0] _GEN_507 = 9'h7 == rs2[8:0] ? coeffs_7 : _GEN_506;
  wire [31:0] _GEN_508 = 9'h8 == rs2[8:0] ? coeffs_8 : _GEN_507;
  wire [31:0] _GEN_509 = 9'h9 == rs2[8:0] ? coeffs_9 : _GEN_508;
  wire [31:0] _GEN_510 = 9'ha == rs2[8:0] ? coeffs_10 : _GEN_509;
  wire [31:0] _GEN_511 = 9'hb == rs2[8:0] ? coeffs_11 : _GEN_510;
  wire [31:0] _GEN_512 = 9'hc == rs2[8:0] ? coeffs_12 : _GEN_511;
  wire [31:0] _GEN_513 = 9'hd == rs2[8:0] ? coeffs_13 : _GEN_512;
  wire [31:0] _GEN_514 = 9'he == rs2[8:0] ? coeffs_14 : _GEN_513;
  wire [31:0] _GEN_515 = 9'hf == rs2[8:0] ? coeffs_15 : _GEN_514;
  wire [31:0] _GEN_516 = 9'h10 == rs2[8:0] ? coeffs_16 : _GEN_515;
  wire [31:0] _GEN_517 = 9'h11 == rs2[8:0] ? coeffs_17 : _GEN_516;
  wire [31:0] _GEN_518 = 9'h12 == rs2[8:0] ? coeffs_18 : _GEN_517;
  wire [31:0] _GEN_519 = 9'h13 == rs2[8:0] ? coeffs_19 : _GEN_518;
  wire [31:0] _GEN_520 = 9'h14 == rs2[8:0] ? coeffs_20 : _GEN_519;
  wire [31:0] _GEN_521 = 9'h15 == rs2[8:0] ? coeffs_21 : _GEN_520;
  wire [31:0] _GEN_522 = 9'h16 == rs2[8:0] ? coeffs_22 : _GEN_521;
  wire [31:0] _GEN_523 = 9'h17 == rs2[8:0] ? coeffs_23 : _GEN_522;
  wire [31:0] _GEN_524 = 9'h18 == rs2[8:0] ? coeffs_24 : _GEN_523;
  wire [31:0] _GEN_525 = 9'h19 == rs2[8:0] ? coeffs_25 : _GEN_524;
  wire [31:0] _GEN_526 = 9'h1a == rs2[8:0] ? coeffs_26 : _GEN_525;
  wire [31:0] _GEN_527 = 9'h1b == rs2[8:0] ? coeffs_27 : _GEN_526;
  wire [31:0] _GEN_528 = 9'h1c == rs2[8:0] ? coeffs_28 : _GEN_527;
  wire [31:0] _GEN_529 = 9'h1d == rs2[8:0] ? coeffs_29 : _GEN_528;
  wire [31:0] _GEN_530 = 9'h1e == rs2[8:0] ? coeffs_30 : _GEN_529;
  wire [31:0] _GEN_531 = 9'h1f == rs2[8:0] ? coeffs_31 : _GEN_530;
  wire [31:0] _GEN_532 = 9'h20 == rs2[8:0] ? coeffs_32 : _GEN_531;
  wire [31:0] _GEN_533 = 9'h21 == rs2[8:0] ? coeffs_33 : _GEN_532;
  wire [31:0] _GEN_534 = 9'h22 == rs2[8:0] ? coeffs_34 : _GEN_533;
  wire [31:0] _GEN_535 = 9'h23 == rs2[8:0] ? coeffs_35 : _GEN_534;
  wire [31:0] _GEN_536 = 9'h24 == rs2[8:0] ? coeffs_36 : _GEN_535;
  wire [31:0] _GEN_537 = 9'h25 == rs2[8:0] ? coeffs_37 : _GEN_536;
  wire [31:0] _GEN_538 = 9'h26 == rs2[8:0] ? coeffs_38 : _GEN_537;
  wire [31:0] _GEN_539 = 9'h27 == rs2[8:0] ? coeffs_39 : _GEN_538;
  wire [31:0] _GEN_540 = 9'h28 == rs2[8:0] ? coeffs_40 : _GEN_539;
  wire [31:0] _GEN_541 = 9'h29 == rs2[8:0] ? coeffs_41 : _GEN_540;
  wire [31:0] _GEN_542 = 9'h2a == rs2[8:0] ? coeffs_42 : _GEN_541;
  wire [31:0] _GEN_543 = 9'h2b == rs2[8:0] ? coeffs_43 : _GEN_542;
  wire [31:0] _GEN_544 = 9'h2c == rs2[8:0] ? coeffs_44 : _GEN_543;
  wire [31:0] _GEN_545 = 9'h2d == rs2[8:0] ? coeffs_45 : _GEN_544;
  wire [31:0] _GEN_546 = 9'h2e == rs2[8:0] ? coeffs_46 : _GEN_545;
  wire [31:0] _GEN_547 = 9'h2f == rs2[8:0] ? coeffs_47 : _GEN_546;
  wire [31:0] _GEN_548 = 9'h30 == rs2[8:0] ? coeffs_48 : _GEN_547;
  wire [31:0] _GEN_549 = 9'h31 == rs2[8:0] ? coeffs_49 : _GEN_548;
  wire [31:0] _GEN_550 = 9'h32 == rs2[8:0] ? coeffs_50 : _GEN_549;
  wire [31:0] _GEN_551 = 9'h33 == rs2[8:0] ? coeffs_51 : _GEN_550;
  wire [31:0] _GEN_552 = 9'h34 == rs2[8:0] ? coeffs_52 : _GEN_551;
  wire [31:0] _GEN_553 = 9'h35 == rs2[8:0] ? coeffs_53 : _GEN_552;
  wire [31:0] _GEN_554 = 9'h36 == rs2[8:0] ? coeffs_54 : _GEN_553;
  wire [31:0] _GEN_555 = 9'h37 == rs2[8:0] ? coeffs_55 : _GEN_554;
  wire [31:0] _GEN_556 = 9'h38 == rs2[8:0] ? coeffs_56 : _GEN_555;
  wire [31:0] _GEN_557 = 9'h39 == rs2[8:0] ? coeffs_57 : _GEN_556;
  wire [31:0] _GEN_558 = 9'h3a == rs2[8:0] ? coeffs_58 : _GEN_557;
  wire [31:0] _GEN_559 = 9'h3b == rs2[8:0] ? coeffs_59 : _GEN_558;
  wire [31:0] _GEN_560 = 9'h3c == rs2[8:0] ? coeffs_60 : _GEN_559;
  wire [31:0] _GEN_561 = 9'h3d == rs2[8:0] ? coeffs_61 : _GEN_560;
  wire [31:0] _GEN_562 = 9'h3e == rs2[8:0] ? coeffs_62 : _GEN_561;
  wire [31:0] _GEN_563 = 9'h3f == rs2[8:0] ? coeffs_63 : _GEN_562;
  wire [31:0] _GEN_564 = 9'h40 == rs2[8:0] ? coeffs_64 : _GEN_563;
  wire [31:0] _GEN_565 = 9'h41 == rs2[8:0] ? coeffs_65 : _GEN_564;
  wire [31:0] _GEN_566 = 9'h42 == rs2[8:0] ? coeffs_66 : _GEN_565;
  wire [31:0] _GEN_567 = 9'h43 == rs2[8:0] ? coeffs_67 : _GEN_566;
  wire [31:0] _GEN_568 = 9'h44 == rs2[8:0] ? coeffs_68 : _GEN_567;
  wire [31:0] _GEN_569 = 9'h45 == rs2[8:0] ? coeffs_69 : _GEN_568;
  wire [31:0] _GEN_570 = 9'h46 == rs2[8:0] ? coeffs_70 : _GEN_569;
  wire [31:0] _GEN_571 = 9'h47 == rs2[8:0] ? coeffs_71 : _GEN_570;
  wire [31:0] _GEN_572 = 9'h48 == rs2[8:0] ? coeffs_72 : _GEN_571;
  wire [31:0] _GEN_573 = 9'h49 == rs2[8:0] ? coeffs_73 : _GEN_572;
  wire [31:0] _GEN_574 = 9'h4a == rs2[8:0] ? coeffs_74 : _GEN_573;
  wire [31:0] _GEN_575 = 9'h4b == rs2[8:0] ? coeffs_75 : _GEN_574;
  wire [31:0] _GEN_576 = 9'h4c == rs2[8:0] ? coeffs_76 : _GEN_575;
  wire [31:0] _GEN_577 = 9'h4d == rs2[8:0] ? coeffs_77 : _GEN_576;
  wire [31:0] _GEN_578 = 9'h4e == rs2[8:0] ? coeffs_78 : _GEN_577;
  wire [31:0] _GEN_579 = 9'h4f == rs2[8:0] ? coeffs_79 : _GEN_578;
  wire [31:0] _GEN_580 = 9'h50 == rs2[8:0] ? coeffs_80 : _GEN_579;
  wire [31:0] _GEN_581 = 9'h51 == rs2[8:0] ? coeffs_81 : _GEN_580;
  wire [31:0] _GEN_582 = 9'h52 == rs2[8:0] ? coeffs_82 : _GEN_581;
  wire [31:0] _GEN_583 = 9'h53 == rs2[8:0] ? coeffs_83 : _GEN_582;
  wire [31:0] _GEN_584 = 9'h54 == rs2[8:0] ? coeffs_84 : _GEN_583;
  wire [31:0] _GEN_585 = 9'h55 == rs2[8:0] ? coeffs_85 : _GEN_584;
  wire [31:0] _GEN_586 = 9'h56 == rs2[8:0] ? coeffs_86 : _GEN_585;
  wire [31:0] _GEN_587 = 9'h57 == rs2[8:0] ? coeffs_87 : _GEN_586;
  wire [31:0] _GEN_588 = 9'h58 == rs2[8:0] ? coeffs_88 : _GEN_587;
  wire [31:0] _GEN_589 = 9'h59 == rs2[8:0] ? coeffs_89 : _GEN_588;
  wire [31:0] _GEN_590 = 9'h5a == rs2[8:0] ? coeffs_90 : _GEN_589;
  wire [31:0] _GEN_591 = 9'h5b == rs2[8:0] ? coeffs_91 : _GEN_590;
  wire [31:0] _GEN_592 = 9'h5c == rs2[8:0] ? coeffs_92 : _GEN_591;
  wire [31:0] _GEN_593 = 9'h5d == rs2[8:0] ? coeffs_93 : _GEN_592;
  wire [31:0] _GEN_594 = 9'h5e == rs2[8:0] ? coeffs_94 : _GEN_593;
  wire [31:0] _GEN_595 = 9'h5f == rs2[8:0] ? coeffs_95 : _GEN_594;
  wire [31:0] _GEN_596 = 9'h60 == rs2[8:0] ? coeffs_96 : _GEN_595;
  wire [31:0] _GEN_597 = 9'h61 == rs2[8:0] ? coeffs_97 : _GEN_596;
  wire [31:0] _GEN_598 = 9'h62 == rs2[8:0] ? coeffs_98 : _GEN_597;
  wire [31:0] _GEN_599 = 9'h63 == rs2[8:0] ? coeffs_99 : _GEN_598;
  wire [31:0] _GEN_600 = 9'h64 == rs2[8:0] ? coeffs_100 : _GEN_599;
  wire [31:0] _GEN_601 = 9'h65 == rs2[8:0] ? coeffs_101 : _GEN_600;
  wire [31:0] _GEN_602 = 9'h66 == rs2[8:0] ? coeffs_102 : _GEN_601;
  wire [31:0] _GEN_603 = 9'h67 == rs2[8:0] ? coeffs_103 : _GEN_602;
  wire [31:0] _GEN_604 = 9'h68 == rs2[8:0] ? coeffs_104 : _GEN_603;
  wire [31:0] _GEN_605 = 9'h69 == rs2[8:0] ? coeffs_105 : _GEN_604;
  wire [31:0] _GEN_606 = 9'h6a == rs2[8:0] ? coeffs_106 : _GEN_605;
  wire [31:0] _GEN_607 = 9'h6b == rs2[8:0] ? coeffs_107 : _GEN_606;
  wire [31:0] _GEN_608 = 9'h6c == rs2[8:0] ? coeffs_108 : _GEN_607;
  wire [31:0] _GEN_609 = 9'h6d == rs2[8:0] ? coeffs_109 : _GEN_608;
  wire [31:0] _GEN_610 = 9'h6e == rs2[8:0] ? coeffs_110 : _GEN_609;
  wire [31:0] _GEN_611 = 9'h6f == rs2[8:0] ? coeffs_111 : _GEN_610;
  wire [31:0] _GEN_612 = 9'h70 == rs2[8:0] ? coeffs_112 : _GEN_611;
  wire [31:0] _GEN_613 = 9'h71 == rs2[8:0] ? coeffs_113 : _GEN_612;
  wire [31:0] _GEN_614 = 9'h72 == rs2[8:0] ? coeffs_114 : _GEN_613;
  wire [31:0] _GEN_615 = 9'h73 == rs2[8:0] ? coeffs_115 : _GEN_614;
  wire [31:0] _GEN_616 = 9'h74 == rs2[8:0] ? coeffs_116 : _GEN_615;
  wire [31:0] _GEN_617 = 9'h75 == rs2[8:0] ? coeffs_117 : _GEN_616;
  wire [31:0] _GEN_618 = 9'h76 == rs2[8:0] ? coeffs_118 : _GEN_617;
  wire [31:0] _GEN_619 = 9'h77 == rs2[8:0] ? coeffs_119 : _GEN_618;
  wire [31:0] _GEN_620 = 9'h78 == rs2[8:0] ? coeffs_120 : _GEN_619;
  wire [31:0] _GEN_621 = 9'h79 == rs2[8:0] ? coeffs_121 : _GEN_620;
  wire [31:0] _GEN_622 = 9'h7a == rs2[8:0] ? coeffs_122 : _GEN_621;
  wire [31:0] _GEN_623 = 9'h7b == rs2[8:0] ? coeffs_123 : _GEN_622;
  wire [31:0] _GEN_624 = 9'h7c == rs2[8:0] ? coeffs_124 : _GEN_623;
  wire [31:0] _GEN_625 = 9'h7d == rs2[8:0] ? coeffs_125 : _GEN_624;
  wire [31:0] _GEN_626 = 9'h7e == rs2[8:0] ? coeffs_126 : _GEN_625;
  wire [31:0] _GEN_627 = 9'h7f == rs2[8:0] ? coeffs_127 : _GEN_626;
  wire [31:0] _GEN_628 = 9'h80 == rs2[8:0] ? coeffs_128 : _GEN_627;
  wire [31:0] _GEN_629 = 9'h81 == rs2[8:0] ? coeffs_129 : _GEN_628;
  wire [31:0] _GEN_630 = 9'h82 == rs2[8:0] ? coeffs_130 : _GEN_629;
  wire [31:0] _GEN_631 = 9'h83 == rs2[8:0] ? coeffs_131 : _GEN_630;
  wire [31:0] _GEN_632 = 9'h84 == rs2[8:0] ? coeffs_132 : _GEN_631;
  wire [31:0] _GEN_633 = 9'h85 == rs2[8:0] ? coeffs_133 : _GEN_632;
  wire [31:0] _GEN_634 = 9'h86 == rs2[8:0] ? coeffs_134 : _GEN_633;
  wire [31:0] _GEN_635 = 9'h87 == rs2[8:0] ? coeffs_135 : _GEN_634;
  wire [31:0] _GEN_636 = 9'h88 == rs2[8:0] ? coeffs_136 : _GEN_635;
  wire [31:0] _GEN_637 = 9'h89 == rs2[8:0] ? coeffs_137 : _GEN_636;
  wire [31:0] _GEN_638 = 9'h8a == rs2[8:0] ? coeffs_138 : _GEN_637;
  wire [31:0] _GEN_639 = 9'h8b == rs2[8:0] ? coeffs_139 : _GEN_638;
  wire [31:0] _GEN_640 = 9'h8c == rs2[8:0] ? coeffs_140 : _GEN_639;
  wire [31:0] _GEN_641 = 9'h8d == rs2[8:0] ? coeffs_141 : _GEN_640;
  wire [31:0] _GEN_642 = 9'h8e == rs2[8:0] ? coeffs_142 : _GEN_641;
  wire [31:0] _GEN_643 = 9'h8f == rs2[8:0] ? coeffs_143 : _GEN_642;
  wire [31:0] _GEN_644 = 9'h90 == rs2[8:0] ? coeffs_144 : _GEN_643;
  wire [31:0] _GEN_645 = 9'h91 == rs2[8:0] ? coeffs_145 : _GEN_644;
  wire [31:0] _GEN_646 = 9'h92 == rs2[8:0] ? coeffs_146 : _GEN_645;
  wire [31:0] _GEN_647 = 9'h93 == rs2[8:0] ? coeffs_147 : _GEN_646;
  wire [31:0] _GEN_648 = 9'h94 == rs2[8:0] ? coeffs_148 : _GEN_647;
  wire [31:0] _GEN_649 = 9'h95 == rs2[8:0] ? coeffs_149 : _GEN_648;
  wire [31:0] _GEN_650 = 9'h96 == rs2[8:0] ? coeffs_150 : _GEN_649;
  wire [31:0] _GEN_651 = 9'h97 == rs2[8:0] ? coeffs_151 : _GEN_650;
  wire [31:0] _GEN_652 = 9'h98 == rs2[8:0] ? coeffs_152 : _GEN_651;
  wire [31:0] _GEN_653 = 9'h99 == rs2[8:0] ? coeffs_153 : _GEN_652;
  wire [31:0] _GEN_654 = 9'h9a == rs2[8:0] ? coeffs_154 : _GEN_653;
  wire [31:0] _GEN_655 = 9'h9b == rs2[8:0] ? coeffs_155 : _GEN_654;
  wire [31:0] _GEN_656 = 9'h9c == rs2[8:0] ? coeffs_156 : _GEN_655;
  wire [31:0] _GEN_657 = 9'h9d == rs2[8:0] ? coeffs_157 : _GEN_656;
  wire [31:0] _GEN_658 = 9'h9e == rs2[8:0] ? coeffs_158 : _GEN_657;
  wire [31:0] _GEN_659 = 9'h9f == rs2[8:0] ? coeffs_159 : _GEN_658;
  wire [31:0] _GEN_660 = 9'ha0 == rs2[8:0] ? coeffs_160 : _GEN_659;
  wire [31:0] _GEN_661 = 9'ha1 == rs2[8:0] ? coeffs_161 : _GEN_660;
  wire [31:0] _GEN_662 = 9'ha2 == rs2[8:0] ? coeffs_162 : _GEN_661;
  wire [31:0] _GEN_663 = 9'ha3 == rs2[8:0] ? coeffs_163 : _GEN_662;
  wire [31:0] _GEN_664 = 9'ha4 == rs2[8:0] ? coeffs_164 : _GEN_663;
  wire [31:0] _GEN_665 = 9'ha5 == rs2[8:0] ? coeffs_165 : _GEN_664;
  wire [31:0] _GEN_666 = 9'ha6 == rs2[8:0] ? coeffs_166 : _GEN_665;
  wire [31:0] _GEN_667 = 9'ha7 == rs2[8:0] ? coeffs_167 : _GEN_666;
  wire [31:0] _GEN_668 = 9'ha8 == rs2[8:0] ? coeffs_168 : _GEN_667;
  wire [31:0] _GEN_669 = 9'ha9 == rs2[8:0] ? coeffs_169 : _GEN_668;
  wire [31:0] _GEN_670 = 9'haa == rs2[8:0] ? coeffs_170 : _GEN_669;
  wire [31:0] _GEN_671 = 9'hab == rs2[8:0] ? coeffs_171 : _GEN_670;
  wire [31:0] _GEN_672 = 9'hac == rs2[8:0] ? coeffs_172 : _GEN_671;
  wire [31:0] _GEN_673 = 9'had == rs2[8:0] ? coeffs_173 : _GEN_672;
  wire [31:0] _GEN_674 = 9'hae == rs2[8:0] ? coeffs_174 : _GEN_673;
  wire [31:0] _GEN_675 = 9'haf == rs2[8:0] ? coeffs_175 : _GEN_674;
  wire [31:0] _GEN_676 = 9'hb0 == rs2[8:0] ? coeffs_176 : _GEN_675;
  wire [31:0] _GEN_677 = 9'hb1 == rs2[8:0] ? coeffs_177 : _GEN_676;
  wire [31:0] _GEN_678 = 9'hb2 == rs2[8:0] ? coeffs_178 : _GEN_677;
  wire [31:0] _GEN_679 = 9'hb3 == rs2[8:0] ? coeffs_179 : _GEN_678;
  wire [31:0] _GEN_680 = 9'hb4 == rs2[8:0] ? coeffs_180 : _GEN_679;
  wire [31:0] _GEN_681 = 9'hb5 == rs2[8:0] ? coeffs_181 : _GEN_680;
  wire [31:0] _GEN_682 = 9'hb6 == rs2[8:0] ? coeffs_182 : _GEN_681;
  wire [31:0] _GEN_683 = 9'hb7 == rs2[8:0] ? coeffs_183 : _GEN_682;
  wire [31:0] _GEN_684 = 9'hb8 == rs2[8:0] ? coeffs_184 : _GEN_683;
  wire [31:0] _GEN_685 = 9'hb9 == rs2[8:0] ? coeffs_185 : _GEN_684;
  wire [31:0] _GEN_686 = 9'hba == rs2[8:0] ? coeffs_186 : _GEN_685;
  wire [31:0] _GEN_687 = 9'hbb == rs2[8:0] ? coeffs_187 : _GEN_686;
  wire [31:0] _GEN_688 = 9'hbc == rs2[8:0] ? coeffs_188 : _GEN_687;
  wire [31:0] _GEN_689 = 9'hbd == rs2[8:0] ? coeffs_189 : _GEN_688;
  wire [31:0] _GEN_690 = 9'hbe == rs2[8:0] ? coeffs_190 : _GEN_689;
  wire [31:0] _GEN_691 = 9'hbf == rs2[8:0] ? coeffs_191 : _GEN_690;
  wire [31:0] _GEN_692 = 9'hc0 == rs2[8:0] ? coeffs_192 : _GEN_691;
  wire [31:0] _GEN_693 = 9'hc1 == rs2[8:0] ? coeffs_193 : _GEN_692;
  wire [31:0] _GEN_694 = 9'hc2 == rs2[8:0] ? coeffs_194 : _GEN_693;
  wire [31:0] _GEN_695 = 9'hc3 == rs2[8:0] ? coeffs_195 : _GEN_694;
  wire [31:0] _GEN_696 = 9'hc4 == rs2[8:0] ? coeffs_196 : _GEN_695;
  wire [31:0] _GEN_697 = 9'hc5 == rs2[8:0] ? coeffs_197 : _GEN_696;
  wire [31:0] _GEN_698 = 9'hc6 == rs2[8:0] ? coeffs_198 : _GEN_697;
  wire [31:0] _GEN_699 = 9'hc7 == rs2[8:0] ? coeffs_199 : _GEN_698;
  wire [31:0] _GEN_700 = 9'hc8 == rs2[8:0] ? coeffs_200 : _GEN_699;
  wire [31:0] _GEN_701 = 9'hc9 == rs2[8:0] ? coeffs_201 : _GEN_700;
  wire [31:0] _GEN_702 = 9'hca == rs2[8:0] ? coeffs_202 : _GEN_701;
  wire [31:0] _GEN_703 = 9'hcb == rs2[8:0] ? coeffs_203 : _GEN_702;
  wire [31:0] _GEN_704 = 9'hcc == rs2[8:0] ? coeffs_204 : _GEN_703;
  wire [31:0] _GEN_705 = 9'hcd == rs2[8:0] ? coeffs_205 : _GEN_704;
  wire [31:0] _GEN_706 = 9'hce == rs2[8:0] ? coeffs_206 : _GEN_705;
  wire [31:0] _GEN_707 = 9'hcf == rs2[8:0] ? coeffs_207 : _GEN_706;
  wire [31:0] _GEN_708 = 9'hd0 == rs2[8:0] ? coeffs_208 : _GEN_707;
  wire [31:0] _GEN_709 = 9'hd1 == rs2[8:0] ? coeffs_209 : _GEN_708;
  wire [31:0] _GEN_710 = 9'hd2 == rs2[8:0] ? coeffs_210 : _GEN_709;
  wire [31:0] _GEN_711 = 9'hd3 == rs2[8:0] ? coeffs_211 : _GEN_710;
  wire [31:0] _GEN_712 = 9'hd4 == rs2[8:0] ? coeffs_212 : _GEN_711;
  wire [31:0] _GEN_713 = 9'hd5 == rs2[8:0] ? coeffs_213 : _GEN_712;
  wire [31:0] _GEN_714 = 9'hd6 == rs2[8:0] ? coeffs_214 : _GEN_713;
  wire [31:0] _GEN_715 = 9'hd7 == rs2[8:0] ? coeffs_215 : _GEN_714;
  wire [31:0] _GEN_716 = 9'hd8 == rs2[8:0] ? coeffs_216 : _GEN_715;
  wire [31:0] _GEN_717 = 9'hd9 == rs2[8:0] ? coeffs_217 : _GEN_716;
  wire [31:0] _GEN_718 = 9'hda == rs2[8:0] ? coeffs_218 : _GEN_717;
  wire [31:0] _GEN_719 = 9'hdb == rs2[8:0] ? coeffs_219 : _GEN_718;
  wire [31:0] _GEN_720 = 9'hdc == rs2[8:0] ? coeffs_220 : _GEN_719;
  wire [31:0] _GEN_721 = 9'hdd == rs2[8:0] ? coeffs_221 : _GEN_720;
  wire [31:0] _GEN_722 = 9'hde == rs2[8:0] ? coeffs_222 : _GEN_721;
  wire [31:0] _GEN_723 = 9'hdf == rs2[8:0] ? coeffs_223 : _GEN_722;
  wire [31:0] _GEN_724 = 9'he0 == rs2[8:0] ? coeffs_224 : _GEN_723;
  wire [31:0] _GEN_725 = 9'he1 == rs2[8:0] ? coeffs_225 : _GEN_724;
  wire [31:0] _GEN_726 = 9'he2 == rs2[8:0] ? coeffs_226 : _GEN_725;
  wire [31:0] _GEN_727 = 9'he3 == rs2[8:0] ? coeffs_227 : _GEN_726;
  wire [31:0] _GEN_728 = 9'he4 == rs2[8:0] ? coeffs_228 : _GEN_727;
  wire [31:0] _GEN_729 = 9'he5 == rs2[8:0] ? coeffs_229 : _GEN_728;
  wire [31:0] _GEN_730 = 9'he6 == rs2[8:0] ? coeffs_230 : _GEN_729;
  wire [31:0] _GEN_731 = 9'he7 == rs2[8:0] ? coeffs_231 : _GEN_730;
  wire [31:0] _GEN_732 = 9'he8 == rs2[8:0] ? coeffs_232 : _GEN_731;
  wire [31:0] _GEN_733 = 9'he9 == rs2[8:0] ? coeffs_233 : _GEN_732;
  wire [31:0] _GEN_734 = 9'hea == rs2[8:0] ? coeffs_234 : _GEN_733;
  wire [31:0] _GEN_735 = 9'heb == rs2[8:0] ? coeffs_235 : _GEN_734;
  wire [31:0] _GEN_736 = 9'hec == rs2[8:0] ? coeffs_236 : _GEN_735;
  wire [31:0] _GEN_737 = 9'hed == rs2[8:0] ? coeffs_237 : _GEN_736;
  wire [31:0] _GEN_738 = 9'hee == rs2[8:0] ? coeffs_238 : _GEN_737;
  wire [31:0] _GEN_739 = 9'hef == rs2[8:0] ? coeffs_239 : _GEN_738;
  wire [31:0] _GEN_740 = 9'hf0 == rs2[8:0] ? coeffs_240 : _GEN_739;
  wire [31:0] _GEN_741 = 9'hf1 == rs2[8:0] ? coeffs_241 : _GEN_740;
  wire [31:0] _GEN_742 = 9'hf2 == rs2[8:0] ? coeffs_242 : _GEN_741;
  wire [31:0] _GEN_743 = 9'hf3 == rs2[8:0] ? coeffs_243 : _GEN_742;
  wire [31:0] _GEN_744 = 9'hf4 == rs2[8:0] ? coeffs_244 : _GEN_743;
  wire [31:0] _GEN_745 = 9'hf5 == rs2[8:0] ? coeffs_245 : _GEN_744;
  wire [31:0] _GEN_746 = 9'hf6 == rs2[8:0] ? coeffs_246 : _GEN_745;
  wire [31:0] _GEN_747 = 9'hf7 == rs2[8:0] ? coeffs_247 : _GEN_746;
  wire [31:0] _GEN_748 = 9'hf8 == rs2[8:0] ? coeffs_248 : _GEN_747;
  wire [31:0] _GEN_749 = 9'hf9 == rs2[8:0] ? coeffs_249 : _GEN_748;
  wire [31:0] _GEN_750 = 9'hfa == rs2[8:0] ? coeffs_250 : _GEN_749;
  wire [31:0] _GEN_751 = 9'hfb == rs2[8:0] ? coeffs_251 : _GEN_750;
  wire [31:0] _GEN_752 = 9'hfc == rs2[8:0] ? coeffs_252 : _GEN_751;
  wire [31:0] _GEN_753 = 9'hfd == rs2[8:0] ? coeffs_253 : _GEN_752;
  wire [31:0] _GEN_754 = 9'hfe == rs2[8:0] ? coeffs_254 : _GEN_753;
  wire [31:0] _GEN_755 = 9'hff == rs2[8:0] ? coeffs_255 : _GEN_754;
  wire [31:0] _GEN_756 = 9'h100 == rs2[8:0] ? coeffs_256 : _GEN_755;
  wire [31:0] _GEN_757 = 9'h101 == rs2[8:0] ? coeffs_257 : _GEN_756;
  wire [31:0] _GEN_758 = 9'h102 == rs2[8:0] ? coeffs_258 : _GEN_757;
  wire [31:0] _GEN_759 = 9'h103 == rs2[8:0] ? coeffs_259 : _GEN_758;
  wire [31:0] _GEN_760 = 9'h104 == rs2[8:0] ? coeffs_260 : _GEN_759;
  wire [31:0] _GEN_761 = 9'h105 == rs2[8:0] ? coeffs_261 : _GEN_760;
  wire [31:0] _GEN_762 = 9'h106 == rs2[8:0] ? coeffs_262 : _GEN_761;
  wire [31:0] _GEN_763 = 9'h107 == rs2[8:0] ? coeffs_263 : _GEN_762;
  wire [31:0] _GEN_764 = 9'h108 == rs2[8:0] ? coeffs_264 : _GEN_763;
  wire [31:0] _GEN_765 = 9'h109 == rs2[8:0] ? coeffs_265 : _GEN_764;
  wire [31:0] _GEN_766 = 9'h10a == rs2[8:0] ? coeffs_266 : _GEN_765;
  wire [31:0] _GEN_767 = 9'h10b == rs2[8:0] ? coeffs_267 : _GEN_766;
  wire [31:0] _GEN_768 = 9'h10c == rs2[8:0] ? coeffs_268 : _GEN_767;
  wire [31:0] _GEN_769 = 9'h10d == rs2[8:0] ? coeffs_269 : _GEN_768;
  wire [31:0] _GEN_770 = 9'h10e == rs2[8:0] ? coeffs_270 : _GEN_769;
  wire [31:0] _GEN_771 = 9'h10f == rs2[8:0] ? coeffs_271 : _GEN_770;
  wire [31:0] _GEN_772 = 9'h110 == rs2[8:0] ? coeffs_272 : _GEN_771;
  wire [31:0] _GEN_773 = 9'h111 == rs2[8:0] ? coeffs_273 : _GEN_772;
  wire [31:0] _GEN_774 = 9'h112 == rs2[8:0] ? coeffs_274 : _GEN_773;
  wire [31:0] _GEN_775 = 9'h113 == rs2[8:0] ? coeffs_275 : _GEN_774;
  wire [31:0] _GEN_776 = 9'h114 == rs2[8:0] ? coeffs_276 : _GEN_775;
  wire [31:0] _GEN_777 = 9'h115 == rs2[8:0] ? coeffs_277 : _GEN_776;
  wire [31:0] _GEN_778 = 9'h116 == rs2[8:0] ? coeffs_278 : _GEN_777;
  wire [31:0] _GEN_779 = 9'h117 == rs2[8:0] ? coeffs_279 : _GEN_778;
  wire [31:0] _GEN_780 = 9'h118 == rs2[8:0] ? coeffs_280 : _GEN_779;
  wire [31:0] _GEN_781 = 9'h119 == rs2[8:0] ? coeffs_281 : _GEN_780;
  wire [31:0] _GEN_782 = 9'h11a == rs2[8:0] ? coeffs_282 : _GEN_781;
  wire [31:0] _GEN_783 = 9'h11b == rs2[8:0] ? coeffs_283 : _GEN_782;
  wire [31:0] _GEN_784 = 9'h11c == rs2[8:0] ? coeffs_284 : _GEN_783;
  wire [31:0] _GEN_785 = 9'h11d == rs2[8:0] ? coeffs_285 : _GEN_784;
  wire [31:0] _GEN_786 = 9'h11e == rs2[8:0] ? coeffs_286 : _GEN_785;
  wire [31:0] _GEN_787 = 9'h11f == rs2[8:0] ? coeffs_287 : _GEN_786;
  wire [31:0] _GEN_788 = 9'h120 == rs2[8:0] ? coeffs_288 : _GEN_787;
  wire [31:0] _GEN_789 = 9'h121 == rs2[8:0] ? coeffs_289 : _GEN_788;
  wire [31:0] _GEN_790 = 9'h122 == rs2[8:0] ? coeffs_290 : _GEN_789;
  wire [31:0] _GEN_791 = 9'h123 == rs2[8:0] ? coeffs_291 : _GEN_790;
  wire [31:0] _GEN_792 = 9'h124 == rs2[8:0] ? coeffs_292 : _GEN_791;
  wire [31:0] _GEN_793 = 9'h125 == rs2[8:0] ? coeffs_293 : _GEN_792;
  wire [31:0] _GEN_794 = 9'h126 == rs2[8:0] ? coeffs_294 : _GEN_793;
  wire [31:0] _GEN_795 = 9'h127 == rs2[8:0] ? coeffs_295 : _GEN_794;
  wire [31:0] _GEN_796 = 9'h128 == rs2[8:0] ? coeffs_296 : _GEN_795;
  wire [31:0] _GEN_797 = 9'h129 == rs2[8:0] ? coeffs_297 : _GEN_796;
  wire [31:0] _GEN_798 = 9'h12a == rs2[8:0] ? coeffs_298 : _GEN_797;
  wire [31:0] _GEN_799 = 9'h12b == rs2[8:0] ? coeffs_299 : _GEN_798;
  wire [31:0] _GEN_800 = 9'h12c == rs2[8:0] ? coeffs_300 : _GEN_799;
  wire [31:0] _GEN_801 = 9'h12d == rs2[8:0] ? coeffs_301 : _GEN_800;
  wire [31:0] _GEN_802 = 9'h12e == rs2[8:0] ? coeffs_302 : _GEN_801;
  wire [31:0] _GEN_803 = 9'h12f == rs2[8:0] ? coeffs_303 : _GEN_802;
  wire [31:0] _GEN_804 = 9'h130 == rs2[8:0] ? coeffs_304 : _GEN_803;
  wire [31:0] _GEN_805 = 9'h131 == rs2[8:0] ? coeffs_305 : _GEN_804;
  wire [31:0] _GEN_806 = 9'h132 == rs2[8:0] ? coeffs_306 : _GEN_805;
  wire [31:0] _GEN_807 = 9'h133 == rs2[8:0] ? coeffs_307 : _GEN_806;
  wire [31:0] _GEN_808 = 9'h134 == rs2[8:0] ? coeffs_308 : _GEN_807;
  wire [31:0] _GEN_809 = 9'h135 == rs2[8:0] ? coeffs_309 : _GEN_808;
  wire [31:0] _GEN_810 = 9'h136 == rs2[8:0] ? coeffs_310 : _GEN_809;
  wire [31:0] _GEN_811 = 9'h137 == rs2[8:0] ? coeffs_311 : _GEN_810;
  wire [31:0] _GEN_812 = 9'h138 == rs2[8:0] ? coeffs_312 : _GEN_811;
  wire [31:0] _GEN_813 = 9'h139 == rs2[8:0] ? coeffs_313 : _GEN_812;
  wire [31:0] _GEN_814 = 9'h13a == rs2[8:0] ? coeffs_314 : _GEN_813;
  wire [31:0] _GEN_815 = 9'h13b == rs2[8:0] ? coeffs_315 : _GEN_814;
  wire [31:0] _GEN_816 = 9'h13c == rs2[8:0] ? coeffs_316 : _GEN_815;
  wire [31:0] _GEN_817 = 9'h13d == rs2[8:0] ? coeffs_317 : _GEN_816;
  wire [31:0] _GEN_818 = 9'h13e == rs2[8:0] ? coeffs_318 : _GEN_817;
  wire [31:0] _GEN_819 = 9'h13f == rs2[8:0] ? coeffs_319 : _GEN_818;
  wire [31:0] _GEN_820 = 9'h140 == rs2[8:0] ? coeffs_320 : _GEN_819;
  wire [31:0] _GEN_821 = 9'h141 == rs2[8:0] ? coeffs_321 : _GEN_820;
  wire [31:0] _GEN_822 = 9'h142 == rs2[8:0] ? coeffs_322 : _GEN_821;
  wire [31:0] _GEN_823 = 9'h143 == rs2[8:0] ? coeffs_323 : _GEN_822;
  wire [31:0] _GEN_824 = 9'h144 == rs2[8:0] ? coeffs_324 : _GEN_823;
  wire [31:0] _GEN_825 = 9'h145 == rs2[8:0] ? coeffs_325 : _GEN_824;
  wire [31:0] _GEN_826 = 9'h146 == rs2[8:0] ? coeffs_326 : _GEN_825;
  wire [31:0] _GEN_827 = 9'h147 == rs2[8:0] ? coeffs_327 : _GEN_826;
  wire [31:0] _GEN_828 = 9'h148 == rs2[8:0] ? coeffs_328 : _GEN_827;
  wire [31:0] _GEN_829 = 9'h149 == rs2[8:0] ? coeffs_329 : _GEN_828;
  wire [31:0] _GEN_830 = 9'h14a == rs2[8:0] ? coeffs_330 : _GEN_829;
  wire [31:0] _GEN_831 = 9'h14b == rs2[8:0] ? coeffs_331 : _GEN_830;
  wire [31:0] _GEN_832 = 9'h14c == rs2[8:0] ? coeffs_332 : _GEN_831;
  wire [31:0] _GEN_833 = 9'h14d == rs2[8:0] ? coeffs_333 : _GEN_832;
  wire [31:0] _GEN_834 = 9'h14e == rs2[8:0] ? coeffs_334 : _GEN_833;
  wire [31:0] _GEN_835 = 9'h14f == rs2[8:0] ? coeffs_335 : _GEN_834;
  wire [31:0] _GEN_836 = 9'h150 == rs2[8:0] ? coeffs_336 : _GEN_835;
  wire [31:0] _GEN_837 = 9'h151 == rs2[8:0] ? coeffs_337 : _GEN_836;
  wire [31:0] _GEN_838 = 9'h152 == rs2[8:0] ? coeffs_338 : _GEN_837;
  wire [31:0] _GEN_839 = 9'h153 == rs2[8:0] ? coeffs_339 : _GEN_838;
  wire [31:0] _GEN_840 = 9'h154 == rs2[8:0] ? coeffs_340 : _GEN_839;
  wire [31:0] _GEN_841 = 9'h155 == rs2[8:0] ? coeffs_341 : _GEN_840;
  wire [31:0] _GEN_842 = 9'h156 == rs2[8:0] ? coeffs_342 : _GEN_841;
  wire [31:0] _GEN_843 = 9'h157 == rs2[8:0] ? coeffs_343 : _GEN_842;
  wire [31:0] _GEN_844 = 9'h158 == rs2[8:0] ? coeffs_344 : _GEN_843;
  wire [31:0] _GEN_845 = 9'h159 == rs2[8:0] ? coeffs_345 : _GEN_844;
  wire [31:0] _GEN_846 = 9'h15a == rs2[8:0] ? coeffs_346 : _GEN_845;
  wire [31:0] _GEN_847 = 9'h15b == rs2[8:0] ? coeffs_347 : _GEN_846;
  wire [31:0] _GEN_848 = 9'h15c == rs2[8:0] ? coeffs_348 : _GEN_847;
  wire [31:0] _GEN_849 = 9'h15d == rs2[8:0] ? coeffs_349 : _GEN_848;
  wire [31:0] _GEN_850 = 9'h15e == rs2[8:0] ? coeffs_350 : _GEN_849;
  wire [31:0] _GEN_851 = 9'h15f == rs2[8:0] ? coeffs_351 : _GEN_850;
  wire [31:0] _GEN_852 = 9'h160 == rs2[8:0] ? coeffs_352 : _GEN_851;
  wire [31:0] _GEN_853 = 9'h161 == rs2[8:0] ? coeffs_353 : _GEN_852;
  wire [31:0] _GEN_854 = 9'h162 == rs2[8:0] ? coeffs_354 : _GEN_853;
  wire [31:0] _GEN_855 = 9'h163 == rs2[8:0] ? coeffs_355 : _GEN_854;
  wire [31:0] _GEN_856 = 9'h164 == rs2[8:0] ? coeffs_356 : _GEN_855;
  wire [31:0] _GEN_857 = 9'h165 == rs2[8:0] ? coeffs_357 : _GEN_856;
  wire [31:0] _GEN_858 = 9'h166 == rs2[8:0] ? coeffs_358 : _GEN_857;
  wire [31:0] _GEN_859 = 9'h167 == rs2[8:0] ? coeffs_359 : _GEN_858;
  wire [31:0] _GEN_860 = 9'h168 == rs2[8:0] ? coeffs_360 : _GEN_859;
  wire [31:0] _GEN_861 = 9'h169 == rs2[8:0] ? coeffs_361 : _GEN_860;
  wire [31:0] _GEN_862 = 9'h16a == rs2[8:0] ? coeffs_362 : _GEN_861;
  wire [31:0] _GEN_863 = 9'h16b == rs2[8:0] ? coeffs_363 : _GEN_862;
  wire [31:0] _GEN_864 = 9'h16c == rs2[8:0] ? coeffs_364 : _GEN_863;
  wire [31:0] _GEN_865 = 9'h16d == rs2[8:0] ? coeffs_365 : _GEN_864;
  wire [31:0] _GEN_866 = 9'h16e == rs2[8:0] ? coeffs_366 : _GEN_865;
  wire [31:0] _GEN_867 = 9'h16f == rs2[8:0] ? coeffs_367 : _GEN_866;
  wire [31:0] _GEN_868 = 9'h170 == rs2[8:0] ? coeffs_368 : _GEN_867;
  wire [31:0] _GEN_869 = 9'h171 == rs2[8:0] ? coeffs_369 : _GEN_868;
  wire [31:0] _GEN_870 = 9'h172 == rs2[8:0] ? coeffs_370 : _GEN_869;
  wire [31:0] _GEN_871 = 9'h173 == rs2[8:0] ? coeffs_371 : _GEN_870;
  wire [31:0] _GEN_872 = 9'h174 == rs2[8:0] ? coeffs_372 : _GEN_871;
  wire [31:0] _GEN_873 = 9'h175 == rs2[8:0] ? coeffs_373 : _GEN_872;
  wire [31:0] _GEN_874 = 9'h176 == rs2[8:0] ? coeffs_374 : _GEN_873;
  wire [31:0] _GEN_875 = 9'h177 == rs2[8:0] ? coeffs_375 : _GEN_874;
  wire [31:0] _GEN_876 = 9'h178 == rs2[8:0] ? coeffs_376 : _GEN_875;
  wire [31:0] _GEN_877 = 9'h179 == rs2[8:0] ? coeffs_377 : _GEN_876;
  wire [31:0] _GEN_878 = 9'h17a == rs2[8:0] ? coeffs_378 : _GEN_877;
  wire [31:0] _GEN_879 = 9'h17b == rs2[8:0] ? coeffs_379 : _GEN_878;
  wire [31:0] _GEN_880 = 9'h17c == rs2[8:0] ? coeffs_380 : _GEN_879;
  wire [31:0] _GEN_881 = 9'h17d == rs2[8:0] ? coeffs_381 : _GEN_880;
  wire [31:0] _GEN_882 = 9'h17e == rs2[8:0] ? coeffs_382 : _GEN_881;
  wire [31:0] _GEN_883 = 9'h17f == rs2[8:0] ? coeffs_383 : _GEN_882;
  wire [31:0] _GEN_884 = 9'h180 == rs2[8:0] ? coeffs_384 : _GEN_883;
  wire [31:0] _GEN_885 = 9'h181 == rs2[8:0] ? coeffs_385 : _GEN_884;
  wire [31:0] _GEN_886 = 9'h182 == rs2[8:0] ? coeffs_386 : _GEN_885;
  wire [31:0] _GEN_887 = 9'h183 == rs2[8:0] ? coeffs_387 : _GEN_886;
  wire [31:0] _GEN_888 = 9'h184 == rs2[8:0] ? coeffs_388 : _GEN_887;
  wire [31:0] _GEN_889 = 9'h185 == rs2[8:0] ? coeffs_389 : _GEN_888;
  wire [31:0] _GEN_890 = 9'h186 == rs2[8:0] ? coeffs_390 : _GEN_889;
  wire [31:0] _GEN_891 = 9'h187 == rs2[8:0] ? coeffs_391 : _GEN_890;
  wire [31:0] _GEN_892 = 9'h188 == rs2[8:0] ? coeffs_392 : _GEN_891;
  wire [31:0] _GEN_893 = 9'h189 == rs2[8:0] ? coeffs_393 : _GEN_892;
  wire [31:0] _GEN_894 = 9'h18a == rs2[8:0] ? coeffs_394 : _GEN_893;
  wire [31:0] _GEN_895 = 9'h18b == rs2[8:0] ? coeffs_395 : _GEN_894;
  wire [31:0] _GEN_896 = 9'h18c == rs2[8:0] ? coeffs_396 : _GEN_895;
  wire [31:0] _GEN_897 = 9'h18d == rs2[8:0] ? coeffs_397 : _GEN_896;
  wire [31:0] _GEN_898 = 9'h18e == rs2[8:0] ? coeffs_398 : _GEN_897;
  wire [31:0] _GEN_899 = 9'h18f == rs2[8:0] ? coeffs_399 : _GEN_898;
  wire [31:0] _GEN_900 = 9'h190 == rs2[8:0] ? coeffs_400 : _GEN_899;
  wire [31:0] _GEN_901 = 9'h191 == rs2[8:0] ? coeffs_401 : _GEN_900;
  wire [31:0] _GEN_902 = 9'h192 == rs2[8:0] ? coeffs_402 : _GEN_901;
  wire [31:0] _GEN_903 = 9'h193 == rs2[8:0] ? coeffs_403 : _GEN_902;
  wire [31:0] _GEN_904 = 9'h194 == rs2[8:0] ? coeffs_404 : _GEN_903;
  wire [31:0] _GEN_905 = 9'h195 == rs2[8:0] ? coeffs_405 : _GEN_904;
  wire [31:0] _GEN_906 = 9'h196 == rs2[8:0] ? coeffs_406 : _GEN_905;
  wire [31:0] _GEN_907 = 9'h197 == rs2[8:0] ? coeffs_407 : _GEN_906;
  wire [31:0] _GEN_908 = 9'h198 == rs2[8:0] ? coeffs_408 : _GEN_907;
  wire [31:0] _GEN_909 = 9'h199 == rs2[8:0] ? coeffs_409 : _GEN_908;
  wire [31:0] _GEN_910 = 9'h19a == rs2[8:0] ? coeffs_410 : _GEN_909;
  wire [31:0] _GEN_911 = 9'h19b == rs2[8:0] ? coeffs_411 : _GEN_910;
  wire [31:0] _GEN_912 = 9'h19c == rs2[8:0] ? coeffs_412 : _GEN_911;
  wire [31:0] _GEN_913 = 9'h19d == rs2[8:0] ? coeffs_413 : _GEN_912;
  wire [31:0] _GEN_914 = 9'h19e == rs2[8:0] ? coeffs_414 : _GEN_913;
  wire [31:0] _GEN_915 = 9'h19f == rs2[8:0] ? coeffs_415 : _GEN_914;
  wire [31:0] _GEN_916 = 9'h1a0 == rs2[8:0] ? coeffs_416 : _GEN_915;
  wire [31:0] _GEN_917 = 9'h1a1 == rs2[8:0] ? coeffs_417 : _GEN_916;
  wire [31:0] _GEN_918 = 9'h1a2 == rs2[8:0] ? coeffs_418 : _GEN_917;
  wire [31:0] _GEN_919 = 9'h1a3 == rs2[8:0] ? coeffs_419 : _GEN_918;
  wire [31:0] _GEN_920 = 9'h1a4 == rs2[8:0] ? coeffs_420 : _GEN_919;
  wire [31:0] _GEN_921 = 9'h1a5 == rs2[8:0] ? coeffs_421 : _GEN_920;
  wire [31:0] _GEN_922 = 9'h1a6 == rs2[8:0] ? coeffs_422 : _GEN_921;
  wire [31:0] _GEN_923 = 9'h1a7 == rs2[8:0] ? coeffs_423 : _GEN_922;
  wire [31:0] _GEN_924 = 9'h1a8 == rs2[8:0] ? coeffs_424 : _GEN_923;
  wire [31:0] _GEN_925 = 9'h1a9 == rs2[8:0] ? coeffs_425 : _GEN_924;
  wire [31:0] _GEN_926 = 9'h1aa == rs2[8:0] ? coeffs_426 : _GEN_925;
  wire [31:0] _GEN_927 = 9'h1ab == rs2[8:0] ? coeffs_427 : _GEN_926;
  wire [31:0] _GEN_928 = 9'h1ac == rs2[8:0] ? coeffs_428 : _GEN_927;
  wire [31:0] _GEN_929 = 9'h1ad == rs2[8:0] ? coeffs_429 : _GEN_928;
  wire [31:0] _GEN_930 = 9'h1ae == rs2[8:0] ? coeffs_430 : _GEN_929;
  wire [31:0] _GEN_931 = 9'h1af == rs2[8:0] ? coeffs_431 : _GEN_930;
  wire [31:0] _GEN_932 = 9'h1b0 == rs2[8:0] ? coeffs_432 : _GEN_931;
  wire [31:0] _GEN_933 = 9'h1b1 == rs2[8:0] ? coeffs_433 : _GEN_932;
  wire [31:0] _GEN_934 = 9'h1b2 == rs2[8:0] ? coeffs_434 : _GEN_933;
  wire [31:0] _GEN_935 = 9'h1b3 == rs2[8:0] ? coeffs_435 : _GEN_934;
  wire [31:0] _GEN_936 = 9'h1b4 == rs2[8:0] ? coeffs_436 : _GEN_935;
  wire [31:0] _GEN_937 = 9'h1b5 == rs2[8:0] ? coeffs_437 : _GEN_936;
  wire [31:0] _GEN_938 = 9'h1b6 == rs2[8:0] ? coeffs_438 : _GEN_937;
  wire [31:0] _GEN_939 = 9'h1b7 == rs2[8:0] ? coeffs_439 : _GEN_938;
  wire [31:0] _GEN_940 = 9'h1b8 == rs2[8:0] ? coeffs_440 : _GEN_939;
  wire [31:0] _GEN_941 = 9'h1b9 == rs2[8:0] ? coeffs_441 : _GEN_940;
  wire [31:0] _GEN_942 = 9'h1ba == rs2[8:0] ? coeffs_442 : _GEN_941;
  wire [31:0] _GEN_943 = 9'h1bb == rs2[8:0] ? coeffs_443 : _GEN_942;
  wire [31:0] _GEN_944 = 9'h1bc == rs2[8:0] ? coeffs_444 : _GEN_943;
  wire [31:0] _GEN_945 = 9'h1bd == rs2[8:0] ? coeffs_445 : _GEN_944;
  wire [31:0] _GEN_946 = 9'h1be == rs2[8:0] ? coeffs_446 : _GEN_945;
  wire [31:0] _GEN_947 = 9'h1bf == rs2[8:0] ? coeffs_447 : _GEN_946;
  wire [31:0] _GEN_948 = 9'h1c0 == rs2[8:0] ? coeffs_448 : _GEN_947;
  wire [31:0] _GEN_949 = 9'h1c1 == rs2[8:0] ? coeffs_449 : _GEN_948;
  wire [31:0] _GEN_950 = 9'h1c2 == rs2[8:0] ? coeffs_450 : _GEN_949;
  wire [31:0] _GEN_951 = 9'h1c3 == rs2[8:0] ? coeffs_451 : _GEN_950;
  wire [31:0] _GEN_952 = 9'h1c4 == rs2[8:0] ? coeffs_452 : _GEN_951;
  wire [31:0] _GEN_953 = 9'h1c5 == rs2[8:0] ? coeffs_453 : _GEN_952;
  wire [31:0] _GEN_954 = 9'h1c6 == rs2[8:0] ? coeffs_454 : _GEN_953;
  wire [31:0] _GEN_955 = 9'h1c7 == rs2[8:0] ? coeffs_455 : _GEN_954;
  wire [31:0] _GEN_956 = 9'h1c8 == rs2[8:0] ? coeffs_456 : _GEN_955;
  wire [31:0] _GEN_957 = 9'h1c9 == rs2[8:0] ? coeffs_457 : _GEN_956;
  wire [31:0] _GEN_958 = 9'h1ca == rs2[8:0] ? coeffs_458 : _GEN_957;
  wire [31:0] _GEN_959 = 9'h1cb == rs2[8:0] ? coeffs_459 : _GEN_958;
  wire [31:0] _GEN_960 = 9'h1cc == rs2[8:0] ? coeffs_460 : _GEN_959;
  wire [31:0] _GEN_961 = 9'h1cd == rs2[8:0] ? coeffs_461 : _GEN_960;
  wire [31:0] _GEN_962 = 9'h1ce == rs2[8:0] ? coeffs_462 : _GEN_961;
  wire [31:0] _GEN_963 = 9'h1cf == rs2[8:0] ? coeffs_463 : _GEN_962;
  wire [31:0] _GEN_964 = 9'h1d0 == rs2[8:0] ? coeffs_464 : _GEN_963;
  wire [31:0] _GEN_965 = 9'h1d1 == rs2[8:0] ? coeffs_465 : _GEN_964;
  wire [31:0] _GEN_966 = 9'h1d2 == rs2[8:0] ? coeffs_466 : _GEN_965;
  wire [31:0] _GEN_967 = 9'h1d3 == rs2[8:0] ? coeffs_467 : _GEN_966;
  wire [31:0] _GEN_968 = 9'h1d4 == rs2[8:0] ? coeffs_468 : _GEN_967;
  wire [31:0] _GEN_969 = 9'h1d5 == rs2[8:0] ? coeffs_469 : _GEN_968;
  wire [31:0] _GEN_970 = 9'h1d6 == rs2[8:0] ? coeffs_470 : _GEN_969;
  wire [31:0] _GEN_971 = 9'h1d7 == rs2[8:0] ? coeffs_471 : _GEN_970;
  wire [31:0] _GEN_972 = 9'h1d8 == rs2[8:0] ? coeffs_472 : _GEN_971;
  wire [31:0] _GEN_973 = 9'h1d9 == rs2[8:0] ? coeffs_473 : _GEN_972;
  wire [31:0] _GEN_974 = 9'h1da == rs2[8:0] ? coeffs_474 : _GEN_973;
  wire [31:0] _GEN_975 = 9'h1db == rs2[8:0] ? coeffs_475 : _GEN_974;
  wire [31:0] _GEN_976 = 9'h1dc == rs2[8:0] ? coeffs_476 : _GEN_975;
  wire [31:0] _GEN_977 = 9'h1dd == rs2[8:0] ? coeffs_477 : _GEN_976;
  wire [31:0] _GEN_978 = 9'h1de == rs2[8:0] ? coeffs_478 : _GEN_977;
  wire [31:0] _GEN_979 = 9'h1df == rs2[8:0] ? coeffs_479 : _GEN_978;
  wire [31:0] _GEN_980 = 9'h1e0 == rs2[8:0] ? coeffs_480 : _GEN_979;
  wire [31:0] _GEN_981 = 9'h1e1 == rs2[8:0] ? coeffs_481 : _GEN_980;
  wire [31:0] _GEN_982 = 9'h1e2 == rs2[8:0] ? coeffs_482 : _GEN_981;
  wire [31:0] _GEN_983 = 9'h1e3 == rs2[8:0] ? coeffs_483 : _GEN_982;
  wire [31:0] _GEN_984 = 9'h1e4 == rs2[8:0] ? coeffs_484 : _GEN_983;
  wire [31:0] _GEN_985 = 9'h1e5 == rs2[8:0] ? coeffs_485 : _GEN_984;
  wire [31:0] _GEN_986 = 9'h1e6 == rs2[8:0] ? coeffs_486 : _GEN_985;
  wire [31:0] _GEN_987 = 9'h1e7 == rs2[8:0] ? coeffs_487 : _GEN_986;
  wire [31:0] _GEN_988 = 9'h1e8 == rs2[8:0] ? coeffs_488 : _GEN_987;
  wire [31:0] _GEN_989 = 9'h1e9 == rs2[8:0] ? coeffs_489 : _GEN_988;
  wire [31:0] _GEN_990 = 9'h1ea == rs2[8:0] ? coeffs_490 : _GEN_989;
  wire [31:0] _GEN_991 = 9'h1eb == rs2[8:0] ? coeffs_491 : _GEN_990;
  wire [31:0] _GEN_992 = 9'h1ec == rs2[8:0] ? coeffs_492 : _GEN_991;
  wire [31:0] _GEN_993 = 9'h1ed == rs2[8:0] ? coeffs_493 : _GEN_992;
  wire [31:0] _GEN_994 = 9'h1ee == rs2[8:0] ? coeffs_494 : _GEN_993;
  wire [31:0] _GEN_995 = 9'h1ef == rs2[8:0] ? coeffs_495 : _GEN_994;
  wire [31:0] _GEN_996 = 9'h1f0 == rs2[8:0] ? coeffs_496 : _GEN_995;
  wire [31:0] _GEN_997 = 9'h1f1 == rs2[8:0] ? coeffs_497 : _GEN_996;
  wire [31:0] _GEN_998 = 9'h1f2 == rs2[8:0] ? coeffs_498 : _GEN_997;
  wire [31:0] _GEN_999 = 9'h1f3 == rs2[8:0] ? coeffs_499 : _GEN_998;
  wire [63:0] _result_T_1 = data_0 * coeffs_0;
  wire [63:0] _result_T_2 = data_1 * coeffs_1;
  wire [63:0] _result_T_3 = data_2 * coeffs_2;
  wire [63:0] _result_T_4 = data_3 * coeffs_3;
  wire [63:0] _result_T_5 = data_4 * coeffs_4;
  wire [63:0] _result_T_6 = data_5 * coeffs_5;
  wire [63:0] _result_T_7 = data_6 * coeffs_6;
  wire [63:0] _result_T_8 = data_7 * coeffs_7;
  wire [63:0] _result_T_9 = data_8 * coeffs_8;
  wire [63:0] _result_T_10 = data_9 * coeffs_9;
  wire [63:0] _result_T_11 = data_10 * coeffs_10;
  wire [63:0] _result_T_12 = data_11 * coeffs_11;
  wire [63:0] _result_T_13 = data_12 * coeffs_12;
  wire [63:0] _result_T_14 = data_13 * coeffs_13;
  wire [63:0] _result_T_15 = data_14 * coeffs_14;
  wire [63:0] _result_T_16 = data_15 * coeffs_15;
  wire [63:0] _result_T_17 = data_16 * coeffs_16;
  wire [63:0] _result_T_18 = data_17 * coeffs_17;
  wire [63:0] _result_T_19 = data_18 * coeffs_18;
  wire [63:0] _result_T_20 = data_19 * coeffs_19;
  wire [63:0] _result_T_21 = data_20 * coeffs_20;
  wire [63:0] _result_T_22 = data_21 * coeffs_21;
  wire [63:0] _result_T_23 = data_22 * coeffs_22;
  wire [63:0] _result_T_24 = data_23 * coeffs_23;
  wire [63:0] _result_T_25 = data_24 * coeffs_24;
  wire [63:0] _result_T_26 = data_25 * coeffs_25;
  wire [63:0] _result_T_27 = data_26 * coeffs_26;
  wire [63:0] _result_T_28 = data_27 * coeffs_27;
  wire [63:0] _result_T_29 = data_28 * coeffs_28;
  wire [63:0] _result_T_30 = data_29 * coeffs_29;
  wire [63:0] _result_T_31 = data_30 * coeffs_30;
  wire [63:0] _result_T_32 = data_31 * coeffs_31;
  wire [63:0] _result_T_33 = data_32 * coeffs_32;
  wire [63:0] _result_T_34 = data_33 * coeffs_33;
  wire [63:0] _result_T_35 = data_34 * coeffs_34;
  wire [63:0] _result_T_36 = data_35 * coeffs_35;
  wire [63:0] _result_T_37 = data_36 * coeffs_36;
  wire [63:0] _result_T_38 = data_37 * coeffs_37;
  wire [63:0] _result_T_39 = data_38 * coeffs_38;
  wire [63:0] _result_T_40 = data_39 * coeffs_39;
  wire [63:0] _result_T_41 = data_40 * coeffs_40;
  wire [63:0] _result_T_42 = data_41 * coeffs_41;
  wire [63:0] _result_T_43 = data_42 * coeffs_42;
  wire [63:0] _result_T_44 = data_43 * coeffs_43;
  wire [63:0] _result_T_45 = data_44 * coeffs_44;
  wire [63:0] _result_T_46 = data_45 * coeffs_45;
  wire [63:0] _result_T_47 = data_46 * coeffs_46;
  wire [63:0] _result_T_48 = data_47 * coeffs_47;
  wire [63:0] _result_T_49 = data_48 * coeffs_48;
  wire [63:0] _result_T_50 = data_49 * coeffs_49;
  wire [63:0] _result_T_51 = data_50 * coeffs_50;
  wire [63:0] _result_T_52 = data_51 * coeffs_51;
  wire [63:0] _result_T_53 = data_52 * coeffs_52;
  wire [63:0] _result_T_54 = data_53 * coeffs_53;
  wire [63:0] _result_T_55 = data_54 * coeffs_54;
  wire [63:0] _result_T_56 = data_55 * coeffs_55;
  wire [63:0] _result_T_57 = data_56 * coeffs_56;
  wire [63:0] _result_T_58 = data_57 * coeffs_57;
  wire [63:0] _result_T_59 = data_58 * coeffs_58;
  wire [63:0] _result_T_60 = data_59 * coeffs_59;
  wire [63:0] _result_T_61 = data_60 * coeffs_60;
  wire [63:0] _result_T_62 = data_61 * coeffs_61;
  wire [63:0] _result_T_63 = data_62 * coeffs_62;
  wire [63:0] _result_T_64 = data_63 * coeffs_63;
  wire [63:0] _result_T_65 = data_64 * coeffs_64;
  wire [63:0] _result_T_66 = data_65 * coeffs_65;
  wire [63:0] _result_T_67 = data_66 * coeffs_66;
  wire [63:0] _result_T_68 = data_67 * coeffs_67;
  wire [63:0] _result_T_69 = data_68 * coeffs_68;
  wire [63:0] _result_T_70 = data_69 * coeffs_69;
  wire [63:0] _result_T_71 = data_70 * coeffs_70;
  wire [63:0] _result_T_72 = data_71 * coeffs_71;
  wire [63:0] _result_T_73 = data_72 * coeffs_72;
  wire [63:0] _result_T_74 = data_73 * coeffs_73;
  wire [63:0] _result_T_75 = data_74 * coeffs_74;
  wire [63:0] _result_T_76 = data_75 * coeffs_75;
  wire [63:0] _result_T_77 = data_76 * coeffs_76;
  wire [63:0] _result_T_78 = data_77 * coeffs_77;
  wire [63:0] _result_T_79 = data_78 * coeffs_78;
  wire [63:0] _result_T_80 = data_79 * coeffs_79;
  wire [63:0] _result_T_81 = data_80 * coeffs_80;
  wire [63:0] _result_T_82 = data_81 * coeffs_81;
  wire [63:0] _result_T_83 = data_82 * coeffs_82;
  wire [63:0] _result_T_84 = data_83 * coeffs_83;
  wire [63:0] _result_T_85 = data_84 * coeffs_84;
  wire [63:0] _result_T_86 = data_85 * coeffs_85;
  wire [63:0] _result_T_87 = data_86 * coeffs_86;
  wire [63:0] _result_T_88 = data_87 * coeffs_87;
  wire [63:0] _result_T_89 = data_88 * coeffs_88;
  wire [63:0] _result_T_90 = data_89 * coeffs_89;
  wire [63:0] _result_T_91 = data_90 * coeffs_90;
  wire [63:0] _result_T_92 = data_91 * coeffs_91;
  wire [63:0] _result_T_93 = data_92 * coeffs_92;
  wire [63:0] _result_T_94 = data_93 * coeffs_93;
  wire [63:0] _result_T_95 = data_94 * coeffs_94;
  wire [63:0] _result_T_96 = data_95 * coeffs_95;
  wire [63:0] _result_T_97 = data_96 * coeffs_96;
  wire [63:0] _result_T_98 = data_97 * coeffs_97;
  wire [63:0] _result_T_99 = data_98 * coeffs_98;
  wire [63:0] _result_T_100 = data_99 * coeffs_99;
  wire [63:0] _result_T_101 = data_100 * coeffs_100;
  wire [63:0] _result_T_102 = data_101 * coeffs_101;
  wire [63:0] _result_T_103 = data_102 * coeffs_102;
  wire [63:0] _result_T_104 = data_103 * coeffs_103;
  wire [63:0] _result_T_105 = data_104 * coeffs_104;
  wire [63:0] _result_T_106 = data_105 * coeffs_105;
  wire [63:0] _result_T_107 = data_106 * coeffs_106;
  wire [63:0] _result_T_108 = data_107 * coeffs_107;
  wire [63:0] _result_T_109 = data_108 * coeffs_108;
  wire [63:0] _result_T_110 = data_109 * coeffs_109;
  wire [63:0] _result_T_111 = data_110 * coeffs_110;
  wire [63:0] _result_T_112 = data_111 * coeffs_111;
  wire [63:0] _result_T_113 = data_112 * coeffs_112;
  wire [63:0] _result_T_114 = data_113 * coeffs_113;
  wire [63:0] _result_T_115 = data_114 * coeffs_114;
  wire [63:0] _result_T_116 = data_115 * coeffs_115;
  wire [63:0] _result_T_117 = data_116 * coeffs_116;
  wire [63:0] _result_T_118 = data_117 * coeffs_117;
  wire [63:0] _result_T_119 = data_118 * coeffs_118;
  wire [63:0] _result_T_120 = data_119 * coeffs_119;
  wire [63:0] _result_T_121 = data_120 * coeffs_120;
  wire [63:0] _result_T_122 = data_121 * coeffs_121;
  wire [63:0] _result_T_123 = data_122 * coeffs_122;
  wire [63:0] _result_T_124 = data_123 * coeffs_123;
  wire [63:0] _result_T_125 = data_124 * coeffs_124;
  wire [63:0] _result_T_126 = data_125 * coeffs_125;
  wire [63:0] _result_T_127 = data_126 * coeffs_126;
  wire [63:0] _result_T_128 = data_127 * coeffs_127;
  wire [63:0] _result_T_129 = data_128 * coeffs_128;
  wire [63:0] _result_T_130 = data_129 * coeffs_129;
  wire [63:0] _result_T_131 = data_130 * coeffs_130;
  wire [63:0] _result_T_132 = data_131 * coeffs_131;
  wire [63:0] _result_T_133 = data_132 * coeffs_132;
  wire [63:0] _result_T_134 = data_133 * coeffs_133;
  wire [63:0] _result_T_135 = data_134 * coeffs_134;
  wire [63:0] _result_T_136 = data_135 * coeffs_135;
  wire [63:0] _result_T_137 = data_136 * coeffs_136;
  wire [63:0] _result_T_138 = data_137 * coeffs_137;
  wire [63:0] _result_T_139 = data_138 * coeffs_138;
  wire [63:0] _result_T_140 = data_139 * coeffs_139;
  wire [63:0] _result_T_141 = data_140 * coeffs_140;
  wire [63:0] _result_T_142 = data_141 * coeffs_141;
  wire [63:0] _result_T_143 = data_142 * coeffs_142;
  wire [63:0] _result_T_144 = data_143 * coeffs_143;
  wire [63:0] _result_T_145 = data_144 * coeffs_144;
  wire [63:0] _result_T_146 = data_145 * coeffs_145;
  wire [63:0] _result_T_147 = data_146 * coeffs_146;
  wire [63:0] _result_T_148 = data_147 * coeffs_147;
  wire [63:0] _result_T_149 = data_148 * coeffs_148;
  wire [63:0] _result_T_150 = data_149 * coeffs_149;
  wire [63:0] _result_T_151 = data_150 * coeffs_150;
  wire [63:0] _result_T_152 = data_151 * coeffs_151;
  wire [63:0] _result_T_153 = data_152 * coeffs_152;
  wire [63:0] _result_T_154 = data_153 * coeffs_153;
  wire [63:0] _result_T_155 = data_154 * coeffs_154;
  wire [63:0] _result_T_156 = data_155 * coeffs_155;
  wire [63:0] _result_T_157 = data_156 * coeffs_156;
  wire [63:0] _result_T_158 = data_157 * coeffs_157;
  wire [63:0] _result_T_159 = data_158 * coeffs_158;
  wire [63:0] _result_T_160 = data_159 * coeffs_159;
  wire [63:0] _result_T_161 = data_160 * coeffs_160;
  wire [63:0] _result_T_162 = data_161 * coeffs_161;
  wire [63:0] _result_T_163 = data_162 * coeffs_162;
  wire [63:0] _result_T_164 = data_163 * coeffs_163;
  wire [63:0] _result_T_165 = data_164 * coeffs_164;
  wire [63:0] _result_T_166 = data_165 * coeffs_165;
  wire [63:0] _result_T_167 = data_166 * coeffs_166;
  wire [63:0] _result_T_168 = data_167 * coeffs_167;
  wire [63:0] _result_T_169 = data_168 * coeffs_168;
  wire [63:0] _result_T_170 = data_169 * coeffs_169;
  wire [63:0] _result_T_171 = data_170 * coeffs_170;
  wire [63:0] _result_T_172 = data_171 * coeffs_171;
  wire [63:0] _result_T_173 = data_172 * coeffs_172;
  wire [63:0] _result_T_174 = data_173 * coeffs_173;
  wire [63:0] _result_T_175 = data_174 * coeffs_174;
  wire [63:0] _result_T_176 = data_175 * coeffs_175;
  wire [63:0] _result_T_177 = data_176 * coeffs_176;
  wire [63:0] _result_T_178 = data_177 * coeffs_177;
  wire [63:0] _result_T_179 = data_178 * coeffs_178;
  wire [63:0] _result_T_180 = data_179 * coeffs_179;
  wire [63:0] _result_T_181 = data_180 * coeffs_180;
  wire [63:0] _result_T_182 = data_181 * coeffs_181;
  wire [63:0] _result_T_183 = data_182 * coeffs_182;
  wire [63:0] _result_T_184 = data_183 * coeffs_183;
  wire [63:0] _result_T_185 = data_184 * coeffs_184;
  wire [63:0] _result_T_186 = data_185 * coeffs_185;
  wire [63:0] _result_T_187 = data_186 * coeffs_186;
  wire [63:0] _result_T_188 = data_187 * coeffs_187;
  wire [63:0] _result_T_189 = data_188 * coeffs_188;
  wire [63:0] _result_T_190 = data_189 * coeffs_189;
  wire [63:0] _result_T_191 = data_190 * coeffs_190;
  wire [63:0] _result_T_192 = data_191 * coeffs_191;
  wire [63:0] _result_T_193 = data_192 * coeffs_192;
  wire [63:0] _result_T_194 = data_193 * coeffs_193;
  wire [63:0] _result_T_195 = data_194 * coeffs_194;
  wire [63:0] _result_T_196 = data_195 * coeffs_195;
  wire [63:0] _result_T_197 = data_196 * coeffs_196;
  wire [63:0] _result_T_198 = data_197 * coeffs_197;
  wire [63:0] _result_T_199 = data_198 * coeffs_198;
  wire [63:0] _result_T_200 = data_199 * coeffs_199;
  wire [63:0] _result_T_201 = data_200 * coeffs_200;
  wire [63:0] _result_T_202 = data_201 * coeffs_201;
  wire [63:0] _result_T_203 = data_202 * coeffs_202;
  wire [63:0] _result_T_204 = data_203 * coeffs_203;
  wire [63:0] _result_T_205 = data_204 * coeffs_204;
  wire [63:0] _result_T_206 = data_205 * coeffs_205;
  wire [63:0] _result_T_207 = data_206 * coeffs_206;
  wire [63:0] _result_T_208 = data_207 * coeffs_207;
  wire [63:0] _result_T_209 = data_208 * coeffs_208;
  wire [63:0] _result_T_210 = data_209 * coeffs_209;
  wire [63:0] _result_T_211 = data_210 * coeffs_210;
  wire [63:0] _result_T_212 = data_211 * coeffs_211;
  wire [63:0] _result_T_213 = data_212 * coeffs_212;
  wire [63:0] _result_T_214 = data_213 * coeffs_213;
  wire [63:0] _result_T_215 = data_214 * coeffs_214;
  wire [63:0] _result_T_216 = data_215 * coeffs_215;
  wire [63:0] _result_T_217 = data_216 * coeffs_216;
  wire [63:0] _result_T_218 = data_217 * coeffs_217;
  wire [63:0] _result_T_219 = data_218 * coeffs_218;
  wire [63:0] _result_T_220 = data_219 * coeffs_219;
  wire [63:0] _result_T_221 = data_220 * coeffs_220;
  wire [63:0] _result_T_222 = data_221 * coeffs_221;
  wire [63:0] _result_T_223 = data_222 * coeffs_222;
  wire [63:0] _result_T_224 = data_223 * coeffs_223;
  wire [63:0] _result_T_225 = data_224 * coeffs_224;
  wire [63:0] _result_T_226 = data_225 * coeffs_225;
  wire [63:0] _result_T_227 = data_226 * coeffs_226;
  wire [63:0] _result_T_228 = data_227 * coeffs_227;
  wire [63:0] _result_T_229 = data_228 * coeffs_228;
  wire [63:0] _result_T_230 = data_229 * coeffs_229;
  wire [63:0] _result_T_231 = data_230 * coeffs_230;
  wire [63:0] _result_T_232 = data_231 * coeffs_231;
  wire [63:0] _result_T_233 = data_232 * coeffs_232;
  wire [63:0] _result_T_234 = data_233 * coeffs_233;
  wire [63:0] _result_T_235 = data_234 * coeffs_234;
  wire [63:0] _result_T_236 = data_235 * coeffs_235;
  wire [63:0] _result_T_237 = data_236 * coeffs_236;
  wire [63:0] _result_T_238 = data_237 * coeffs_237;
  wire [63:0] _result_T_239 = data_238 * coeffs_238;
  wire [63:0] _result_T_240 = data_239 * coeffs_239;
  wire [63:0] _result_T_241 = data_240 * coeffs_240;
  wire [63:0] _result_T_242 = data_241 * coeffs_241;
  wire [63:0] _result_T_243 = data_242 * coeffs_242;
  wire [63:0] _result_T_244 = data_243 * coeffs_243;
  wire [63:0] _result_T_245 = data_244 * coeffs_244;
  wire [63:0] _result_T_246 = data_245 * coeffs_245;
  wire [63:0] _result_T_247 = data_246 * coeffs_246;
  wire [63:0] _result_T_248 = data_247 * coeffs_247;
  wire [63:0] _result_T_249 = data_248 * coeffs_248;
  wire [63:0] _result_T_250 = data_249 * coeffs_249;
  wire [63:0] _result_T_251 = data_250 * coeffs_250;
  wire [63:0] _result_T_252 = data_251 * coeffs_251;
  wire [63:0] _result_T_253 = data_252 * coeffs_252;
  wire [63:0] _result_T_254 = data_253 * coeffs_253;
  wire [63:0] _result_T_255 = data_254 * coeffs_254;
  wire [63:0] _result_T_256 = data_255 * coeffs_255;
  wire [63:0] _result_T_257 = data_256 * coeffs_256;
  wire [63:0] _result_T_258 = data_257 * coeffs_257;
  wire [63:0] _result_T_259 = data_258 * coeffs_258;
  wire [63:0] _result_T_260 = data_259 * coeffs_259;
  wire [63:0] _result_T_261 = data_260 * coeffs_260;
  wire [63:0] _result_T_262 = data_261 * coeffs_261;
  wire [63:0] _result_T_263 = data_262 * coeffs_262;
  wire [63:0] _result_T_264 = data_263 * coeffs_263;
  wire [63:0] _result_T_265 = data_264 * coeffs_264;
  wire [63:0] _result_T_266 = data_265 * coeffs_265;
  wire [63:0] _result_T_267 = data_266 * coeffs_266;
  wire [63:0] _result_T_268 = data_267 * coeffs_267;
  wire [63:0] _result_T_269 = data_268 * coeffs_268;
  wire [63:0] _result_T_270 = data_269 * coeffs_269;
  wire [63:0] _result_T_271 = data_270 * coeffs_270;
  wire [63:0] _result_T_272 = data_271 * coeffs_271;
  wire [63:0] _result_T_273 = data_272 * coeffs_272;
  wire [63:0] _result_T_274 = data_273 * coeffs_273;
  wire [63:0] _result_T_275 = data_274 * coeffs_274;
  wire [63:0] _result_T_276 = data_275 * coeffs_275;
  wire [63:0] _result_T_277 = data_276 * coeffs_276;
  wire [63:0] _result_T_278 = data_277 * coeffs_277;
  wire [63:0] _result_T_279 = data_278 * coeffs_278;
  wire [63:0] _result_T_280 = data_279 * coeffs_279;
  wire [63:0] _result_T_281 = data_280 * coeffs_280;
  wire [63:0] _result_T_282 = data_281 * coeffs_281;
  wire [63:0] _result_T_283 = data_282 * coeffs_282;
  wire [63:0] _result_T_284 = data_283 * coeffs_283;
  wire [63:0] _result_T_285 = data_284 * coeffs_284;
  wire [63:0] _result_T_286 = data_285 * coeffs_285;
  wire [63:0] _result_T_287 = data_286 * coeffs_286;
  wire [63:0] _result_T_288 = data_287 * coeffs_287;
  wire [63:0] _result_T_289 = data_288 * coeffs_288;
  wire [63:0] _result_T_290 = data_289 * coeffs_289;
  wire [63:0] _result_T_291 = data_290 * coeffs_290;
  wire [63:0] _result_T_292 = data_291 * coeffs_291;
  wire [63:0] _result_T_293 = data_292 * coeffs_292;
  wire [63:0] _result_T_294 = data_293 * coeffs_293;
  wire [63:0] _result_T_295 = data_294 * coeffs_294;
  wire [63:0] _result_T_296 = data_295 * coeffs_295;
  wire [63:0] _result_T_297 = data_296 * coeffs_296;
  wire [63:0] _result_T_298 = data_297 * coeffs_297;
  wire [63:0] _result_T_299 = data_298 * coeffs_298;
  wire [63:0] _result_T_300 = data_299 * coeffs_299;
  wire [63:0] _result_T_301 = data_300 * coeffs_300;
  wire [63:0] _result_T_302 = data_301 * coeffs_301;
  wire [63:0] _result_T_303 = data_302 * coeffs_302;
  wire [63:0] _result_T_304 = data_303 * coeffs_303;
  wire [63:0] _result_T_305 = data_304 * coeffs_304;
  wire [63:0] _result_T_306 = data_305 * coeffs_305;
  wire [63:0] _result_T_307 = data_306 * coeffs_306;
  wire [63:0] _result_T_308 = data_307 * coeffs_307;
  wire [63:0] _result_T_309 = data_308 * coeffs_308;
  wire [63:0] _result_T_310 = data_309 * coeffs_309;
  wire [63:0] _result_T_311 = data_310 * coeffs_310;
  wire [63:0] _result_T_312 = data_311 * coeffs_311;
  wire [63:0] _result_T_313 = data_312 * coeffs_312;
  wire [63:0] _result_T_314 = data_313 * coeffs_313;
  wire [63:0] _result_T_315 = data_314 * coeffs_314;
  wire [63:0] _result_T_316 = data_315 * coeffs_315;
  wire [63:0] _result_T_317 = data_316 * coeffs_316;
  wire [63:0] _result_T_318 = data_317 * coeffs_317;
  wire [63:0] _result_T_319 = data_318 * coeffs_318;
  wire [63:0] _result_T_320 = data_319 * coeffs_319;
  wire [63:0] _result_T_321 = data_320 * coeffs_320;
  wire [63:0] _result_T_322 = data_321 * coeffs_321;
  wire [63:0] _result_T_323 = data_322 * coeffs_322;
  wire [63:0] _result_T_324 = data_323 * coeffs_323;
  wire [63:0] _result_T_325 = data_324 * coeffs_324;
  wire [63:0] _result_T_326 = data_325 * coeffs_325;
  wire [63:0] _result_T_327 = data_326 * coeffs_326;
  wire [63:0] _result_T_328 = data_327 * coeffs_327;
  wire [63:0] _result_T_329 = data_328 * coeffs_328;
  wire [63:0] _result_T_330 = data_329 * coeffs_329;
  wire [63:0] _result_T_331 = data_330 * coeffs_330;
  wire [63:0] _result_T_332 = data_331 * coeffs_331;
  wire [63:0] _result_T_333 = data_332 * coeffs_332;
  wire [63:0] _result_T_334 = data_333 * coeffs_333;
  wire [63:0] _result_T_335 = data_334 * coeffs_334;
  wire [63:0] _result_T_336 = data_335 * coeffs_335;
  wire [63:0] _result_T_337 = data_336 * coeffs_336;
  wire [63:0] _result_T_338 = data_337 * coeffs_337;
  wire [63:0] _result_T_339 = data_338 * coeffs_338;
  wire [63:0] _result_T_340 = data_339 * coeffs_339;
  wire [63:0] _result_T_341 = data_340 * coeffs_340;
  wire [63:0] _result_T_342 = data_341 * coeffs_341;
  wire [63:0] _result_T_343 = data_342 * coeffs_342;
  wire [63:0] _result_T_344 = data_343 * coeffs_343;
  wire [63:0] _result_T_345 = data_344 * coeffs_344;
  wire [63:0] _result_T_346 = data_345 * coeffs_345;
  wire [63:0] _result_T_347 = data_346 * coeffs_346;
  wire [63:0] _result_T_348 = data_347 * coeffs_347;
  wire [63:0] _result_T_349 = data_348 * coeffs_348;
  wire [63:0] _result_T_350 = data_349 * coeffs_349;
  wire [63:0] _result_T_351 = data_350 * coeffs_350;
  wire [63:0] _result_T_352 = data_351 * coeffs_351;
  wire [63:0] _result_T_353 = data_352 * coeffs_352;
  wire [63:0] _result_T_354 = data_353 * coeffs_353;
  wire [63:0] _result_T_355 = data_354 * coeffs_354;
  wire [63:0] _result_T_356 = data_355 * coeffs_355;
  wire [63:0] _result_T_357 = data_356 * coeffs_356;
  wire [63:0] _result_T_358 = data_357 * coeffs_357;
  wire [63:0] _result_T_359 = data_358 * coeffs_358;
  wire [63:0] _result_T_360 = data_359 * coeffs_359;
  wire [63:0] _result_T_361 = data_360 * coeffs_360;
  wire [63:0] _result_T_362 = data_361 * coeffs_361;
  wire [63:0] _result_T_363 = data_362 * coeffs_362;
  wire [63:0] _result_T_364 = data_363 * coeffs_363;
  wire [63:0] _result_T_365 = data_364 * coeffs_364;
  wire [63:0] _result_T_366 = data_365 * coeffs_365;
  wire [63:0] _result_T_367 = data_366 * coeffs_366;
  wire [63:0] _result_T_368 = data_367 * coeffs_367;
  wire [63:0] _result_T_369 = data_368 * coeffs_368;
  wire [63:0] _result_T_370 = data_369 * coeffs_369;
  wire [63:0] _result_T_371 = data_370 * coeffs_370;
  wire [63:0] _result_T_372 = data_371 * coeffs_371;
  wire [63:0] _result_T_373 = data_372 * coeffs_372;
  wire [63:0] _result_T_374 = data_373 * coeffs_373;
  wire [63:0] _result_T_375 = data_374 * coeffs_374;
  wire [63:0] _result_T_376 = data_375 * coeffs_375;
  wire [63:0] _result_T_377 = data_376 * coeffs_376;
  wire [63:0] _result_T_378 = data_377 * coeffs_377;
  wire [63:0] _result_T_379 = data_378 * coeffs_378;
  wire [63:0] _result_T_380 = data_379 * coeffs_379;
  wire [63:0] _result_T_381 = data_380 * coeffs_380;
  wire [63:0] _result_T_382 = data_381 * coeffs_381;
  wire [63:0] _result_T_383 = data_382 * coeffs_382;
  wire [63:0] _result_T_384 = data_383 * coeffs_383;
  wire [63:0] _result_T_385 = data_384 * coeffs_384;
  wire [63:0] _result_T_386 = data_385 * coeffs_385;
  wire [63:0] _result_T_387 = data_386 * coeffs_386;
  wire [63:0] _result_T_388 = data_387 * coeffs_387;
  wire [63:0] _result_T_389 = data_388 * coeffs_388;
  wire [63:0] _result_T_390 = data_389 * coeffs_389;
  wire [63:0] _result_T_391 = data_390 * coeffs_390;
  wire [63:0] _result_T_392 = data_391 * coeffs_391;
  wire [63:0] _result_T_393 = data_392 * coeffs_392;
  wire [63:0] _result_T_394 = data_393 * coeffs_393;
  wire [63:0] _result_T_395 = data_394 * coeffs_394;
  wire [63:0] _result_T_396 = data_395 * coeffs_395;
  wire [63:0] _result_T_397 = data_396 * coeffs_396;
  wire [63:0] _result_T_398 = data_397 * coeffs_397;
  wire [63:0] _result_T_399 = data_398 * coeffs_398;
  wire [63:0] _result_T_400 = data_399 * coeffs_399;
  wire [63:0] _result_T_401 = data_400 * coeffs_400;
  wire [63:0] _result_T_402 = data_401 * coeffs_401;
  wire [63:0] _result_T_403 = data_402 * coeffs_402;
  wire [63:0] _result_T_404 = data_403 * coeffs_403;
  wire [63:0] _result_T_405 = data_404 * coeffs_404;
  wire [63:0] _result_T_406 = data_405 * coeffs_405;
  wire [63:0] _result_T_407 = data_406 * coeffs_406;
  wire [63:0] _result_T_408 = data_407 * coeffs_407;
  wire [63:0] _result_T_409 = data_408 * coeffs_408;
  wire [63:0] _result_T_410 = data_409 * coeffs_409;
  wire [63:0] _result_T_411 = data_410 * coeffs_410;
  wire [63:0] _result_T_412 = data_411 * coeffs_411;
  wire [63:0] _result_T_413 = data_412 * coeffs_412;
  wire [63:0] _result_T_414 = data_413 * coeffs_413;
  wire [63:0] _result_T_415 = data_414 * coeffs_414;
  wire [63:0] _result_T_416 = data_415 * coeffs_415;
  wire [63:0] _result_T_417 = data_416 * coeffs_416;
  wire [63:0] _result_T_418 = data_417 * coeffs_417;
  wire [63:0] _result_T_419 = data_418 * coeffs_418;
  wire [63:0] _result_T_420 = data_419 * coeffs_419;
  wire [63:0] _result_T_421 = data_420 * coeffs_420;
  wire [63:0] _result_T_422 = data_421 * coeffs_421;
  wire [63:0] _result_T_423 = data_422 * coeffs_422;
  wire [63:0] _result_T_424 = data_423 * coeffs_423;
  wire [63:0] _result_T_425 = data_424 * coeffs_424;
  wire [63:0] _result_T_426 = data_425 * coeffs_425;
  wire [63:0] _result_T_427 = data_426 * coeffs_426;
  wire [63:0] _result_T_428 = data_427 * coeffs_427;
  wire [63:0] _result_T_429 = data_428 * coeffs_428;
  wire [63:0] _result_T_430 = data_429 * coeffs_429;
  wire [63:0] _result_T_431 = data_430 * coeffs_430;
  wire [63:0] _result_T_432 = data_431 * coeffs_431;
  wire [63:0] _result_T_433 = data_432 * coeffs_432;
  wire [63:0] _result_T_434 = data_433 * coeffs_433;
  wire [63:0] _result_T_435 = data_434 * coeffs_434;
  wire [63:0] _result_T_436 = data_435 * coeffs_435;
  wire [63:0] _result_T_437 = data_436 * coeffs_436;
  wire [63:0] _result_T_438 = data_437 * coeffs_437;
  wire [63:0] _result_T_439 = data_438 * coeffs_438;
  wire [63:0] _result_T_440 = data_439 * coeffs_439;
  wire [63:0] _result_T_441 = data_440 * coeffs_440;
  wire [63:0] _result_T_442 = data_441 * coeffs_441;
  wire [63:0] _result_T_443 = data_442 * coeffs_442;
  wire [63:0] _result_T_444 = data_443 * coeffs_443;
  wire [63:0] _result_T_445 = data_444 * coeffs_444;
  wire [63:0] _result_T_446 = data_445 * coeffs_445;
  wire [63:0] _result_T_447 = data_446 * coeffs_446;
  wire [63:0] _result_T_448 = data_447 * coeffs_447;
  wire [63:0] _result_T_449 = data_448 * coeffs_448;
  wire [63:0] _result_T_450 = data_449 * coeffs_449;
  wire [63:0] _result_T_451 = data_450 * coeffs_450;
  wire [63:0] _result_T_452 = data_451 * coeffs_451;
  wire [63:0] _result_T_453 = data_452 * coeffs_452;
  wire [63:0] _result_T_454 = data_453 * coeffs_453;
  wire [63:0] _result_T_455 = data_454 * coeffs_454;
  wire [63:0] _result_T_456 = data_455 * coeffs_455;
  wire [63:0] _result_T_457 = data_456 * coeffs_456;
  wire [63:0] _result_T_458 = data_457 * coeffs_457;
  wire [63:0] _result_T_459 = data_458 * coeffs_458;
  wire [63:0] _result_T_460 = data_459 * coeffs_459;
  wire [63:0] _result_T_461 = data_460 * coeffs_460;
  wire [63:0] _result_T_462 = data_461 * coeffs_461;
  wire [63:0] _result_T_463 = data_462 * coeffs_462;
  wire [63:0] _result_T_464 = data_463 * coeffs_463;
  wire [63:0] _result_T_465 = data_464 * coeffs_464;
  wire [63:0] _result_T_466 = data_465 * coeffs_465;
  wire [63:0] _result_T_467 = data_466 * coeffs_466;
  wire [63:0] _result_T_468 = data_467 * coeffs_467;
  wire [63:0] _result_T_469 = data_468 * coeffs_468;
  wire [63:0] _result_T_470 = data_469 * coeffs_469;
  wire [63:0] _result_T_471 = data_470 * coeffs_470;
  wire [63:0] _result_T_472 = data_471 * coeffs_471;
  wire [63:0] _result_T_473 = data_472 * coeffs_472;
  wire [63:0] _result_T_474 = data_473 * coeffs_473;
  wire [63:0] _result_T_475 = data_474 * coeffs_474;
  wire [63:0] _result_T_476 = data_475 * coeffs_475;
  wire [63:0] _result_T_477 = data_476 * coeffs_476;
  wire [63:0] _result_T_478 = data_477 * coeffs_477;
  wire [63:0] _result_T_479 = data_478 * coeffs_478;
  wire [63:0] _result_T_480 = data_479 * coeffs_479;
  wire [63:0] _result_T_481 = data_480 * coeffs_480;
  wire [63:0] _result_T_482 = data_481 * coeffs_481;
  wire [63:0] _result_T_483 = data_482 * coeffs_482;
  wire [63:0] _result_T_484 = data_483 * coeffs_483;
  wire [63:0] _result_T_485 = data_484 * coeffs_484;
  wire [63:0] _result_T_486 = data_485 * coeffs_485;
  wire [63:0] _result_T_487 = data_486 * coeffs_486;
  wire [63:0] _result_T_488 = data_487 * coeffs_487;
  wire [63:0] _result_T_489 = data_488 * coeffs_488;
  wire [63:0] _result_T_490 = data_489 * coeffs_489;
  wire [63:0] _result_T_491 = data_490 * coeffs_490;
  wire [63:0] _result_T_492 = data_491 * coeffs_491;
  wire [63:0] _result_T_493 = data_492 * coeffs_492;
  wire [63:0] _result_T_494 = data_493 * coeffs_493;
  wire [63:0] _result_T_495 = data_494 * coeffs_494;
  wire [63:0] _result_T_496 = data_495 * coeffs_495;
  wire [63:0] _result_T_497 = data_496 * coeffs_496;
  wire [63:0] _result_T_498 = data_497 * coeffs_497;
  wire [63:0] _result_T_499 = data_498 * coeffs_498;
  wire [63:0] _result_T_500 = data_499 * coeffs_499;
  wire [63:0] _result_T_502 = _result_T_1 + _result_T_2;
  wire [63:0] _result_T_504 = _result_T_502 + _result_T_3;
  wire [63:0] _result_T_506 = _result_T_504 + _result_T_4;
  wire [63:0] _result_T_508 = _result_T_506 + _result_T_5;
  wire [63:0] _result_T_510 = _result_T_508 + _result_T_6;
  wire [63:0] _result_T_512 = _result_T_510 + _result_T_7;
  wire [63:0] _result_T_514 = _result_T_512 + _result_T_8;
  wire [63:0] _result_T_516 = _result_T_514 + _result_T_9;
  wire [63:0] _result_T_518 = _result_T_516 + _result_T_10;
  wire [63:0] _result_T_520 = _result_T_518 + _result_T_11;
  wire [63:0] _result_T_522 = _result_T_520 + _result_T_12;
  wire [63:0] _result_T_524 = _result_T_522 + _result_T_13;
  wire [63:0] _result_T_526 = _result_T_524 + _result_T_14;
  wire [63:0] _result_T_528 = _result_T_526 + _result_T_15;
  wire [63:0] _result_T_530 = _result_T_528 + _result_T_16;
  wire [63:0] _result_T_532 = _result_T_530 + _result_T_17;
  wire [63:0] _result_T_534 = _result_T_532 + _result_T_18;
  wire [63:0] _result_T_536 = _result_T_534 + _result_T_19;
  wire [63:0] _result_T_538 = _result_T_536 + _result_T_20;
  wire [63:0] _result_T_540 = _result_T_538 + _result_T_21;
  wire [63:0] _result_T_542 = _result_T_540 + _result_T_22;
  wire [63:0] _result_T_544 = _result_T_542 + _result_T_23;
  wire [63:0] _result_T_546 = _result_T_544 + _result_T_24;
  wire [63:0] _result_T_548 = _result_T_546 + _result_T_25;
  wire [63:0] _result_T_550 = _result_T_548 + _result_T_26;
  wire [63:0] _result_T_552 = _result_T_550 + _result_T_27;
  wire [63:0] _result_T_554 = _result_T_552 + _result_T_28;
  wire [63:0] _result_T_556 = _result_T_554 + _result_T_29;
  wire [63:0] _result_T_558 = _result_T_556 + _result_T_30;
  wire [63:0] _result_T_560 = _result_T_558 + _result_T_31;
  wire [63:0] _result_T_562 = _result_T_560 + _result_T_32;
  wire [63:0] _result_T_564 = _result_T_562 + _result_T_33;
  wire [63:0] _result_T_566 = _result_T_564 + _result_T_34;
  wire [63:0] _result_T_568 = _result_T_566 + _result_T_35;
  wire [63:0] _result_T_570 = _result_T_568 + _result_T_36;
  wire [63:0] _result_T_572 = _result_T_570 + _result_T_37;
  wire [63:0] _result_T_574 = _result_T_572 + _result_T_38;
  wire [63:0] _result_T_576 = _result_T_574 + _result_T_39;
  wire [63:0] _result_T_578 = _result_T_576 + _result_T_40;
  wire [63:0] _result_T_580 = _result_T_578 + _result_T_41;
  wire [63:0] _result_T_582 = _result_T_580 + _result_T_42;
  wire [63:0] _result_T_584 = _result_T_582 + _result_T_43;
  wire [63:0] _result_T_586 = _result_T_584 + _result_T_44;
  wire [63:0] _result_T_588 = _result_T_586 + _result_T_45;
  wire [63:0] _result_T_590 = _result_T_588 + _result_T_46;
  wire [63:0] _result_T_592 = _result_T_590 + _result_T_47;
  wire [63:0] _result_T_594 = _result_T_592 + _result_T_48;
  wire [63:0] _result_T_596 = _result_T_594 + _result_T_49;
  wire [63:0] _result_T_598 = _result_T_596 + _result_T_50;
  wire [63:0] _result_T_600 = _result_T_598 + _result_T_51;
  wire [63:0] _result_T_602 = _result_T_600 + _result_T_52;
  wire [63:0] _result_T_604 = _result_T_602 + _result_T_53;
  wire [63:0] _result_T_606 = _result_T_604 + _result_T_54;
  wire [63:0] _result_T_608 = _result_T_606 + _result_T_55;
  wire [63:0] _result_T_610 = _result_T_608 + _result_T_56;
  wire [63:0] _result_T_612 = _result_T_610 + _result_T_57;
  wire [63:0] _result_T_614 = _result_T_612 + _result_T_58;
  wire [63:0] _result_T_616 = _result_T_614 + _result_T_59;
  wire [63:0] _result_T_618 = _result_T_616 + _result_T_60;
  wire [63:0] _result_T_620 = _result_T_618 + _result_T_61;
  wire [63:0] _result_T_622 = _result_T_620 + _result_T_62;
  wire [63:0] _result_T_624 = _result_T_622 + _result_T_63;
  wire [63:0] _result_T_626 = _result_T_624 + _result_T_64;
  wire [63:0] _result_T_628 = _result_T_626 + _result_T_65;
  wire [63:0] _result_T_630 = _result_T_628 + _result_T_66;
  wire [63:0] _result_T_632 = _result_T_630 + _result_T_67;
  wire [63:0] _result_T_634 = _result_T_632 + _result_T_68;
  wire [63:0] _result_T_636 = _result_T_634 + _result_T_69;
  wire [63:0] _result_T_638 = _result_T_636 + _result_T_70;
  wire [63:0] _result_T_640 = _result_T_638 + _result_T_71;
  wire [63:0] _result_T_642 = _result_T_640 + _result_T_72;
  wire [63:0] _result_T_644 = _result_T_642 + _result_T_73;
  wire [63:0] _result_T_646 = _result_T_644 + _result_T_74;
  wire [63:0] _result_T_648 = _result_T_646 + _result_T_75;
  wire [63:0] _result_T_650 = _result_T_648 + _result_T_76;
  wire [63:0] _result_T_652 = _result_T_650 + _result_T_77;
  wire [63:0] _result_T_654 = _result_T_652 + _result_T_78;
  wire [63:0] _result_T_656 = _result_T_654 + _result_T_79;
  wire [63:0] _result_T_658 = _result_T_656 + _result_T_80;
  wire [63:0] _result_T_660 = _result_T_658 + _result_T_81;
  wire [63:0] _result_T_662 = _result_T_660 + _result_T_82;
  wire [63:0] _result_T_664 = _result_T_662 + _result_T_83;
  wire [63:0] _result_T_666 = _result_T_664 + _result_T_84;
  wire [63:0] _result_T_668 = _result_T_666 + _result_T_85;
  wire [63:0] _result_T_670 = _result_T_668 + _result_T_86;
  wire [63:0] _result_T_672 = _result_T_670 + _result_T_87;
  wire [63:0] _result_T_674 = _result_T_672 + _result_T_88;
  wire [63:0] _result_T_676 = _result_T_674 + _result_T_89;
  wire [63:0] _result_T_678 = _result_T_676 + _result_T_90;
  wire [63:0] _result_T_680 = _result_T_678 + _result_T_91;
  wire [63:0] _result_T_682 = _result_T_680 + _result_T_92;
  wire [63:0] _result_T_684 = _result_T_682 + _result_T_93;
  wire [63:0] _result_T_686 = _result_T_684 + _result_T_94;
  wire [63:0] _result_T_688 = _result_T_686 + _result_T_95;
  wire [63:0] _result_T_690 = _result_T_688 + _result_T_96;
  wire [63:0] _result_T_692 = _result_T_690 + _result_T_97;
  wire [63:0] _result_T_694 = _result_T_692 + _result_T_98;
  wire [63:0] _result_T_696 = _result_T_694 + _result_T_99;
  wire [63:0] _result_T_698 = _result_T_696 + _result_T_100;
  wire [63:0] _result_T_700 = _result_T_698 + _result_T_101;
  wire [63:0] _result_T_702 = _result_T_700 + _result_T_102;
  wire [63:0] _result_T_704 = _result_T_702 + _result_T_103;
  wire [63:0] _result_T_706 = _result_T_704 + _result_T_104;
  wire [63:0] _result_T_708 = _result_T_706 + _result_T_105;
  wire [63:0] _result_T_710 = _result_T_708 + _result_T_106;
  wire [63:0] _result_T_712 = _result_T_710 + _result_T_107;
  wire [63:0] _result_T_714 = _result_T_712 + _result_T_108;
  wire [63:0] _result_T_716 = _result_T_714 + _result_T_109;
  wire [63:0] _result_T_718 = _result_T_716 + _result_T_110;
  wire [63:0] _result_T_720 = _result_T_718 + _result_T_111;
  wire [63:0] _result_T_722 = _result_T_720 + _result_T_112;
  wire [63:0] _result_T_724 = _result_T_722 + _result_T_113;
  wire [63:0] _result_T_726 = _result_T_724 + _result_T_114;
  wire [63:0] _result_T_728 = _result_T_726 + _result_T_115;
  wire [63:0] _result_T_730 = _result_T_728 + _result_T_116;
  wire [63:0] _result_T_732 = _result_T_730 + _result_T_117;
  wire [63:0] _result_T_734 = _result_T_732 + _result_T_118;
  wire [63:0] _result_T_736 = _result_T_734 + _result_T_119;
  wire [63:0] _result_T_738 = _result_T_736 + _result_T_120;
  wire [63:0] _result_T_740 = _result_T_738 + _result_T_121;
  wire [63:0] _result_T_742 = _result_T_740 + _result_T_122;
  wire [63:0] _result_T_744 = _result_T_742 + _result_T_123;
  wire [63:0] _result_T_746 = _result_T_744 + _result_T_124;
  wire [63:0] _result_T_748 = _result_T_746 + _result_T_125;
  wire [63:0] _result_T_750 = _result_T_748 + _result_T_126;
  wire [63:0] _result_T_752 = _result_T_750 + _result_T_127;
  wire [63:0] _result_T_754 = _result_T_752 + _result_T_128;
  wire [63:0] _result_T_756 = _result_T_754 + _result_T_129;
  wire [63:0] _result_T_758 = _result_T_756 + _result_T_130;
  wire [63:0] _result_T_760 = _result_T_758 + _result_T_131;
  wire [63:0] _result_T_762 = _result_T_760 + _result_T_132;
  wire [63:0] _result_T_764 = _result_T_762 + _result_T_133;
  wire [63:0] _result_T_766 = _result_T_764 + _result_T_134;
  wire [63:0] _result_T_768 = _result_T_766 + _result_T_135;
  wire [63:0] _result_T_770 = _result_T_768 + _result_T_136;
  wire [63:0] _result_T_772 = _result_T_770 + _result_T_137;
  wire [63:0] _result_T_774 = _result_T_772 + _result_T_138;
  wire [63:0] _result_T_776 = _result_T_774 + _result_T_139;
  wire [63:0] _result_T_778 = _result_T_776 + _result_T_140;
  wire [63:0] _result_T_780 = _result_T_778 + _result_T_141;
  wire [63:0] _result_T_782 = _result_T_780 + _result_T_142;
  wire [63:0] _result_T_784 = _result_T_782 + _result_T_143;
  wire [63:0] _result_T_786 = _result_T_784 + _result_T_144;
  wire [63:0] _result_T_788 = _result_T_786 + _result_T_145;
  wire [63:0] _result_T_790 = _result_T_788 + _result_T_146;
  wire [63:0] _result_T_792 = _result_T_790 + _result_T_147;
  wire [63:0] _result_T_794 = _result_T_792 + _result_T_148;
  wire [63:0] _result_T_796 = _result_T_794 + _result_T_149;
  wire [63:0] _result_T_798 = _result_T_796 + _result_T_150;
  wire [63:0] _result_T_800 = _result_T_798 + _result_T_151;
  wire [63:0] _result_T_802 = _result_T_800 + _result_T_152;
  wire [63:0] _result_T_804 = _result_T_802 + _result_T_153;
  wire [63:0] _result_T_806 = _result_T_804 + _result_T_154;
  wire [63:0] _result_T_808 = _result_T_806 + _result_T_155;
  wire [63:0] _result_T_810 = _result_T_808 + _result_T_156;
  wire [63:0] _result_T_812 = _result_T_810 + _result_T_157;
  wire [63:0] _result_T_814 = _result_T_812 + _result_T_158;
  wire [63:0] _result_T_816 = _result_T_814 + _result_T_159;
  wire [63:0] _result_T_818 = _result_T_816 + _result_T_160;
  wire [63:0] _result_T_820 = _result_T_818 + _result_T_161;
  wire [63:0] _result_T_822 = _result_T_820 + _result_T_162;
  wire [63:0] _result_T_824 = _result_T_822 + _result_T_163;
  wire [63:0] _result_T_826 = _result_T_824 + _result_T_164;
  wire [63:0] _result_T_828 = _result_T_826 + _result_T_165;
  wire [63:0] _result_T_830 = _result_T_828 + _result_T_166;
  wire [63:0] _result_T_832 = _result_T_830 + _result_T_167;
  wire [63:0] _result_T_834 = _result_T_832 + _result_T_168;
  wire [63:0] _result_T_836 = _result_T_834 + _result_T_169;
  wire [63:0] _result_T_838 = _result_T_836 + _result_T_170;
  wire [63:0] _result_T_840 = _result_T_838 + _result_T_171;
  wire [63:0] _result_T_842 = _result_T_840 + _result_T_172;
  wire [63:0] _result_T_844 = _result_T_842 + _result_T_173;
  wire [63:0] _result_T_846 = _result_T_844 + _result_T_174;
  wire [63:0] _result_T_848 = _result_T_846 + _result_T_175;
  wire [63:0] _result_T_850 = _result_T_848 + _result_T_176;
  wire [63:0] _result_T_852 = _result_T_850 + _result_T_177;
  wire [63:0] _result_T_854 = _result_T_852 + _result_T_178;
  wire [63:0] _result_T_856 = _result_T_854 + _result_T_179;
  wire [63:0] _result_T_858 = _result_T_856 + _result_T_180;
  wire [63:0] _result_T_860 = _result_T_858 + _result_T_181;
  wire [63:0] _result_T_862 = _result_T_860 + _result_T_182;
  wire [63:0] _result_T_864 = _result_T_862 + _result_T_183;
  wire [63:0] _result_T_866 = _result_T_864 + _result_T_184;
  wire [63:0] _result_T_868 = _result_T_866 + _result_T_185;
  wire [63:0] _result_T_870 = _result_T_868 + _result_T_186;
  wire [63:0] _result_T_872 = _result_T_870 + _result_T_187;
  wire [63:0] _result_T_874 = _result_T_872 + _result_T_188;
  wire [63:0] _result_T_876 = _result_T_874 + _result_T_189;
  wire [63:0] _result_T_878 = _result_T_876 + _result_T_190;
  wire [63:0] _result_T_880 = _result_T_878 + _result_T_191;
  wire [63:0] _result_T_882 = _result_T_880 + _result_T_192;
  wire [63:0] _result_T_884 = _result_T_882 + _result_T_193;
  wire [63:0] _result_T_886 = _result_T_884 + _result_T_194;
  wire [63:0] _result_T_888 = _result_T_886 + _result_T_195;
  wire [63:0] _result_T_890 = _result_T_888 + _result_T_196;
  wire [63:0] _result_T_892 = _result_T_890 + _result_T_197;
  wire [63:0] _result_T_894 = _result_T_892 + _result_T_198;
  wire [63:0] _result_T_896 = _result_T_894 + _result_T_199;
  wire [63:0] _result_T_898 = _result_T_896 + _result_T_200;
  wire [63:0] _result_T_900 = _result_T_898 + _result_T_201;
  wire [63:0] _result_T_902 = _result_T_900 + _result_T_202;
  wire [63:0] _result_T_904 = _result_T_902 + _result_T_203;
  wire [63:0] _result_T_906 = _result_T_904 + _result_T_204;
  wire [63:0] _result_T_908 = _result_T_906 + _result_T_205;
  wire [63:0] _result_T_910 = _result_T_908 + _result_T_206;
  wire [63:0] _result_T_912 = _result_T_910 + _result_T_207;
  wire [63:0] _result_T_914 = _result_T_912 + _result_T_208;
  wire [63:0] _result_T_916 = _result_T_914 + _result_T_209;
  wire [63:0] _result_T_918 = _result_T_916 + _result_T_210;
  wire [63:0] _result_T_920 = _result_T_918 + _result_T_211;
  wire [63:0] _result_T_922 = _result_T_920 + _result_T_212;
  wire [63:0] _result_T_924 = _result_T_922 + _result_T_213;
  wire [63:0] _result_T_926 = _result_T_924 + _result_T_214;
  wire [63:0] _result_T_928 = _result_T_926 + _result_T_215;
  wire [63:0] _result_T_930 = _result_T_928 + _result_T_216;
  wire [63:0] _result_T_932 = _result_T_930 + _result_T_217;
  wire [63:0] _result_T_934 = _result_T_932 + _result_T_218;
  wire [63:0] _result_T_936 = _result_T_934 + _result_T_219;
  wire [63:0] _result_T_938 = _result_T_936 + _result_T_220;
  wire [63:0] _result_T_940 = _result_T_938 + _result_T_221;
  wire [63:0] _result_T_942 = _result_T_940 + _result_T_222;
  wire [63:0] _result_T_944 = _result_T_942 + _result_T_223;
  wire [63:0] _result_T_946 = _result_T_944 + _result_T_224;
  wire [63:0] _result_T_948 = _result_T_946 + _result_T_225;
  wire [63:0] _result_T_950 = _result_T_948 + _result_T_226;
  wire [63:0] _result_T_952 = _result_T_950 + _result_T_227;
  wire [63:0] _result_T_954 = _result_T_952 + _result_T_228;
  wire [63:0] _result_T_956 = _result_T_954 + _result_T_229;
  wire [63:0] _result_T_958 = _result_T_956 + _result_T_230;
  wire [63:0] _result_T_960 = _result_T_958 + _result_T_231;
  wire [63:0] _result_T_962 = _result_T_960 + _result_T_232;
  wire [63:0] _result_T_964 = _result_T_962 + _result_T_233;
  wire [63:0] _result_T_966 = _result_T_964 + _result_T_234;
  wire [63:0] _result_T_968 = _result_T_966 + _result_T_235;
  wire [63:0] _result_T_970 = _result_T_968 + _result_T_236;
  wire [63:0] _result_T_972 = _result_T_970 + _result_T_237;
  wire [63:0] _result_T_974 = _result_T_972 + _result_T_238;
  wire [63:0] _result_T_976 = _result_T_974 + _result_T_239;
  wire [63:0] _result_T_978 = _result_T_976 + _result_T_240;
  wire [63:0] _result_T_980 = _result_T_978 + _result_T_241;
  wire [63:0] _result_T_982 = _result_T_980 + _result_T_242;
  wire [63:0] _result_T_984 = _result_T_982 + _result_T_243;
  wire [63:0] _result_T_986 = _result_T_984 + _result_T_244;
  wire [63:0] _result_T_988 = _result_T_986 + _result_T_245;
  wire [63:0] _result_T_990 = _result_T_988 + _result_T_246;
  wire [63:0] _result_T_992 = _result_T_990 + _result_T_247;
  wire [63:0] _result_T_994 = _result_T_992 + _result_T_248;
  wire [63:0] _result_T_996 = _result_T_994 + _result_T_249;
  wire [63:0] _result_T_998 = _result_T_996 + _result_T_250;
  wire [63:0] _result_T_1000 = _result_T_998 + _result_T_251;
  wire [63:0] _result_T_1002 = _result_T_1000 + _result_T_252;
  wire [63:0] _result_T_1004 = _result_T_1002 + _result_T_253;
  wire [63:0] _result_T_1006 = _result_T_1004 + _result_T_254;
  wire [63:0] _result_T_1008 = _result_T_1006 + _result_T_255;
  wire [63:0] _result_T_1010 = _result_T_1008 + _result_T_256;
  wire [63:0] _result_T_1012 = _result_T_1010 + _result_T_257;
  wire [63:0] _result_T_1014 = _result_T_1012 + _result_T_258;
  wire [63:0] _result_T_1016 = _result_T_1014 + _result_T_259;
  wire [63:0] _result_T_1018 = _result_T_1016 + _result_T_260;
  wire [63:0] _result_T_1020 = _result_T_1018 + _result_T_261;
  wire [63:0] _result_T_1022 = _result_T_1020 + _result_T_262;
  wire [63:0] _result_T_1024 = _result_T_1022 + _result_T_263;
  wire [63:0] _result_T_1026 = _result_T_1024 + _result_T_264;
  wire [63:0] _result_T_1028 = _result_T_1026 + _result_T_265;
  wire [63:0] _result_T_1030 = _result_T_1028 + _result_T_266;
  wire [63:0] _result_T_1032 = _result_T_1030 + _result_T_267;
  wire [63:0] _result_T_1034 = _result_T_1032 + _result_T_268;
  wire [63:0] _result_T_1036 = _result_T_1034 + _result_T_269;
  wire [63:0] _result_T_1038 = _result_T_1036 + _result_T_270;
  wire [63:0] _result_T_1040 = _result_T_1038 + _result_T_271;
  wire [63:0] _result_T_1042 = _result_T_1040 + _result_T_272;
  wire [63:0] _result_T_1044 = _result_T_1042 + _result_T_273;
  wire [63:0] _result_T_1046 = _result_T_1044 + _result_T_274;
  wire [63:0] _result_T_1048 = _result_T_1046 + _result_T_275;
  wire [63:0] _result_T_1050 = _result_T_1048 + _result_T_276;
  wire [63:0] _result_T_1052 = _result_T_1050 + _result_T_277;
  wire [63:0] _result_T_1054 = _result_T_1052 + _result_T_278;
  wire [63:0] _result_T_1056 = _result_T_1054 + _result_T_279;
  wire [63:0] _result_T_1058 = _result_T_1056 + _result_T_280;
  wire [63:0] _result_T_1060 = _result_T_1058 + _result_T_281;
  wire [63:0] _result_T_1062 = _result_T_1060 + _result_T_282;
  wire [63:0] _result_T_1064 = _result_T_1062 + _result_T_283;
  wire [63:0] _result_T_1066 = _result_T_1064 + _result_T_284;
  wire [63:0] _result_T_1068 = _result_T_1066 + _result_T_285;
  wire [63:0] _result_T_1070 = _result_T_1068 + _result_T_286;
  wire [63:0] _result_T_1072 = _result_T_1070 + _result_T_287;
  wire [63:0] _result_T_1074 = _result_T_1072 + _result_T_288;
  wire [63:0] _result_T_1076 = _result_T_1074 + _result_T_289;
  wire [63:0] _result_T_1078 = _result_T_1076 + _result_T_290;
  wire [63:0] _result_T_1080 = _result_T_1078 + _result_T_291;
  wire [63:0] _result_T_1082 = _result_T_1080 + _result_T_292;
  wire [63:0] _result_T_1084 = _result_T_1082 + _result_T_293;
  wire [63:0] _result_T_1086 = _result_T_1084 + _result_T_294;
  wire [63:0] _result_T_1088 = _result_T_1086 + _result_T_295;
  wire [63:0] _result_T_1090 = _result_T_1088 + _result_T_296;
  wire [63:0] _result_T_1092 = _result_T_1090 + _result_T_297;
  wire [63:0] _result_T_1094 = _result_T_1092 + _result_T_298;
  wire [63:0] _result_T_1096 = _result_T_1094 + _result_T_299;
  wire [63:0] _result_T_1098 = _result_T_1096 + _result_T_300;
  wire [63:0] _result_T_1100 = _result_T_1098 + _result_T_301;
  wire [63:0] _result_T_1102 = _result_T_1100 + _result_T_302;
  wire [63:0] _result_T_1104 = _result_T_1102 + _result_T_303;
  wire [63:0] _result_T_1106 = _result_T_1104 + _result_T_304;
  wire [63:0] _result_T_1108 = _result_T_1106 + _result_T_305;
  wire [63:0] _result_T_1110 = _result_T_1108 + _result_T_306;
  wire [63:0] _result_T_1112 = _result_T_1110 + _result_T_307;
  wire [63:0] _result_T_1114 = _result_T_1112 + _result_T_308;
  wire [63:0] _result_T_1116 = _result_T_1114 + _result_T_309;
  wire [63:0] _result_T_1118 = _result_T_1116 + _result_T_310;
  wire [63:0] _result_T_1120 = _result_T_1118 + _result_T_311;
  wire [63:0] _result_T_1122 = _result_T_1120 + _result_T_312;
  wire [63:0] _result_T_1124 = _result_T_1122 + _result_T_313;
  wire [63:0] _result_T_1126 = _result_T_1124 + _result_T_314;
  wire [63:0] _result_T_1128 = _result_T_1126 + _result_T_315;
  wire [63:0] _result_T_1130 = _result_T_1128 + _result_T_316;
  wire [63:0] _result_T_1132 = _result_T_1130 + _result_T_317;
  wire [63:0] _result_T_1134 = _result_T_1132 + _result_T_318;
  wire [63:0] _result_T_1136 = _result_T_1134 + _result_T_319;
  wire [63:0] _result_T_1138 = _result_T_1136 + _result_T_320;
  wire [63:0] _result_T_1140 = _result_T_1138 + _result_T_321;
  wire [63:0] _result_T_1142 = _result_T_1140 + _result_T_322;
  wire [63:0] _result_T_1144 = _result_T_1142 + _result_T_323;
  wire [63:0] _result_T_1146 = _result_T_1144 + _result_T_324;
  wire [63:0] _result_T_1148 = _result_T_1146 + _result_T_325;
  wire [63:0] _result_T_1150 = _result_T_1148 + _result_T_326;
  wire [63:0] _result_T_1152 = _result_T_1150 + _result_T_327;
  wire [63:0] _result_T_1154 = _result_T_1152 + _result_T_328;
  wire [63:0] _result_T_1156 = _result_T_1154 + _result_T_329;
  wire [63:0] _result_T_1158 = _result_T_1156 + _result_T_330;
  wire [63:0] _result_T_1160 = _result_T_1158 + _result_T_331;
  wire [63:0] _result_T_1162 = _result_T_1160 + _result_T_332;
  wire [63:0] _result_T_1164 = _result_T_1162 + _result_T_333;
  wire [63:0] _result_T_1166 = _result_T_1164 + _result_T_334;
  wire [63:0] _result_T_1168 = _result_T_1166 + _result_T_335;
  wire [63:0] _result_T_1170 = _result_T_1168 + _result_T_336;
  wire [63:0] _result_T_1172 = _result_T_1170 + _result_T_337;
  wire [63:0] _result_T_1174 = _result_T_1172 + _result_T_338;
  wire [63:0] _result_T_1176 = _result_T_1174 + _result_T_339;
  wire [63:0] _result_T_1178 = _result_T_1176 + _result_T_340;
  wire [63:0] _result_T_1180 = _result_T_1178 + _result_T_341;
  wire [63:0] _result_T_1182 = _result_T_1180 + _result_T_342;
  wire [63:0] _result_T_1184 = _result_T_1182 + _result_T_343;
  wire [63:0] _result_T_1186 = _result_T_1184 + _result_T_344;
  wire [63:0] _result_T_1188 = _result_T_1186 + _result_T_345;
  wire [63:0] _result_T_1190 = _result_T_1188 + _result_T_346;
  wire [63:0] _result_T_1192 = _result_T_1190 + _result_T_347;
  wire [63:0] _result_T_1194 = _result_T_1192 + _result_T_348;
  wire [63:0] _result_T_1196 = _result_T_1194 + _result_T_349;
  wire [63:0] _result_T_1198 = _result_T_1196 + _result_T_350;
  wire [63:0] _result_T_1200 = _result_T_1198 + _result_T_351;
  wire [63:0] _result_T_1202 = _result_T_1200 + _result_T_352;
  wire [63:0] _result_T_1204 = _result_T_1202 + _result_T_353;
  wire [63:0] _result_T_1206 = _result_T_1204 + _result_T_354;
  wire [63:0] _result_T_1208 = _result_T_1206 + _result_T_355;
  wire [63:0] _result_T_1210 = _result_T_1208 + _result_T_356;
  wire [63:0] _result_T_1212 = _result_T_1210 + _result_T_357;
  wire [63:0] _result_T_1214 = _result_T_1212 + _result_T_358;
  wire [63:0] _result_T_1216 = _result_T_1214 + _result_T_359;
  wire [63:0] _result_T_1218 = _result_T_1216 + _result_T_360;
  wire [63:0] _result_T_1220 = _result_T_1218 + _result_T_361;
  wire [63:0] _result_T_1222 = _result_T_1220 + _result_T_362;
  wire [63:0] _result_T_1224 = _result_T_1222 + _result_T_363;
  wire [63:0] _result_T_1226 = _result_T_1224 + _result_T_364;
  wire [63:0] _result_T_1228 = _result_T_1226 + _result_T_365;
  wire [63:0] _result_T_1230 = _result_T_1228 + _result_T_366;
  wire [63:0] _result_T_1232 = _result_T_1230 + _result_T_367;
  wire [63:0] _result_T_1234 = _result_T_1232 + _result_T_368;
  wire [63:0] _result_T_1236 = _result_T_1234 + _result_T_369;
  wire [63:0] _result_T_1238 = _result_T_1236 + _result_T_370;
  wire [63:0] _result_T_1240 = _result_T_1238 + _result_T_371;
  wire [63:0] _result_T_1242 = _result_T_1240 + _result_T_372;
  wire [63:0] _result_T_1244 = _result_T_1242 + _result_T_373;
  wire [63:0] _result_T_1246 = _result_T_1244 + _result_T_374;
  wire [63:0] _result_T_1248 = _result_T_1246 + _result_T_375;
  wire [63:0] _result_T_1250 = _result_T_1248 + _result_T_376;
  wire [63:0] _result_T_1252 = _result_T_1250 + _result_T_377;
  wire [63:0] _result_T_1254 = _result_T_1252 + _result_T_378;
  wire [63:0] _result_T_1256 = _result_T_1254 + _result_T_379;
  wire [63:0] _result_T_1258 = _result_T_1256 + _result_T_380;
  wire [63:0] _result_T_1260 = _result_T_1258 + _result_T_381;
  wire [63:0] _result_T_1262 = _result_T_1260 + _result_T_382;
  wire [63:0] _result_T_1264 = _result_T_1262 + _result_T_383;
  wire [63:0] _result_T_1266 = _result_T_1264 + _result_T_384;
  wire [63:0] _result_T_1268 = _result_T_1266 + _result_T_385;
  wire [63:0] _result_T_1270 = _result_T_1268 + _result_T_386;
  wire [63:0] _result_T_1272 = _result_T_1270 + _result_T_387;
  wire [63:0] _result_T_1274 = _result_T_1272 + _result_T_388;
  wire [63:0] _result_T_1276 = _result_T_1274 + _result_T_389;
  wire [63:0] _result_T_1278 = _result_T_1276 + _result_T_390;
  wire [63:0] _result_T_1280 = _result_T_1278 + _result_T_391;
  wire [63:0] _result_T_1282 = _result_T_1280 + _result_T_392;
  wire [63:0] _result_T_1284 = _result_T_1282 + _result_T_393;
  wire [63:0] _result_T_1286 = _result_T_1284 + _result_T_394;
  wire [63:0] _result_T_1288 = _result_T_1286 + _result_T_395;
  wire [63:0] _result_T_1290 = _result_T_1288 + _result_T_396;
  wire [63:0] _result_T_1292 = _result_T_1290 + _result_T_397;
  wire [63:0] _result_T_1294 = _result_T_1292 + _result_T_398;
  wire [63:0] _result_T_1296 = _result_T_1294 + _result_T_399;
  wire [63:0] _result_T_1298 = _result_T_1296 + _result_T_400;
  wire [63:0] _result_T_1300 = _result_T_1298 + _result_T_401;
  wire [63:0] _result_T_1302 = _result_T_1300 + _result_T_402;
  wire [63:0] _result_T_1304 = _result_T_1302 + _result_T_403;
  wire [63:0] _result_T_1306 = _result_T_1304 + _result_T_404;
  wire [63:0] _result_T_1308 = _result_T_1306 + _result_T_405;
  wire [63:0] _result_T_1310 = _result_T_1308 + _result_T_406;
  wire [63:0] _result_T_1312 = _result_T_1310 + _result_T_407;
  wire [63:0] _result_T_1314 = _result_T_1312 + _result_T_408;
  wire [63:0] _result_T_1316 = _result_T_1314 + _result_T_409;
  wire [63:0] _result_T_1318 = _result_T_1316 + _result_T_410;
  wire [63:0] _result_T_1320 = _result_T_1318 + _result_T_411;
  wire [63:0] _result_T_1322 = _result_T_1320 + _result_T_412;
  wire [63:0] _result_T_1324 = _result_T_1322 + _result_T_413;
  wire [63:0] _result_T_1326 = _result_T_1324 + _result_T_414;
  wire [63:0] _result_T_1328 = _result_T_1326 + _result_T_415;
  wire [63:0] _result_T_1330 = _result_T_1328 + _result_T_416;
  wire [63:0] _result_T_1332 = _result_T_1330 + _result_T_417;
  wire [63:0] _result_T_1334 = _result_T_1332 + _result_T_418;
  wire [63:0] _result_T_1336 = _result_T_1334 + _result_T_419;
  wire [63:0] _result_T_1338 = _result_T_1336 + _result_T_420;
  wire [63:0] _result_T_1340 = _result_T_1338 + _result_T_421;
  wire [63:0] _result_T_1342 = _result_T_1340 + _result_T_422;
  wire [63:0] _result_T_1344 = _result_T_1342 + _result_T_423;
  wire [63:0] _result_T_1346 = _result_T_1344 + _result_T_424;
  wire [63:0] _result_T_1348 = _result_T_1346 + _result_T_425;
  wire [63:0] _result_T_1350 = _result_T_1348 + _result_T_426;
  wire [63:0] _result_T_1352 = _result_T_1350 + _result_T_427;
  wire [63:0] _result_T_1354 = _result_T_1352 + _result_T_428;
  wire [63:0] _result_T_1356 = _result_T_1354 + _result_T_429;
  wire [63:0] _result_T_1358 = _result_T_1356 + _result_T_430;
  wire [63:0] _result_T_1360 = _result_T_1358 + _result_T_431;
  wire [63:0] _result_T_1362 = _result_T_1360 + _result_T_432;
  wire [63:0] _result_T_1364 = _result_T_1362 + _result_T_433;
  wire [63:0] _result_T_1366 = _result_T_1364 + _result_T_434;
  wire [63:0] _result_T_1368 = _result_T_1366 + _result_T_435;
  wire [63:0] _result_T_1370 = _result_T_1368 + _result_T_436;
  wire [63:0] _result_T_1372 = _result_T_1370 + _result_T_437;
  wire [63:0] _result_T_1374 = _result_T_1372 + _result_T_438;
  wire [63:0] _result_T_1376 = _result_T_1374 + _result_T_439;
  wire [63:0] _result_T_1378 = _result_T_1376 + _result_T_440;
  wire [63:0] _result_T_1380 = _result_T_1378 + _result_T_441;
  wire [63:0] _result_T_1382 = _result_T_1380 + _result_T_442;
  wire [63:0] _result_T_1384 = _result_T_1382 + _result_T_443;
  wire [63:0] _result_T_1386 = _result_T_1384 + _result_T_444;
  wire [63:0] _result_T_1388 = _result_T_1386 + _result_T_445;
  wire [63:0] _result_T_1390 = _result_T_1388 + _result_T_446;
  wire [63:0] _result_T_1392 = _result_T_1390 + _result_T_447;
  wire [63:0] _result_T_1394 = _result_T_1392 + _result_T_448;
  wire [63:0] _result_T_1396 = _result_T_1394 + _result_T_449;
  wire [63:0] _result_T_1398 = _result_T_1396 + _result_T_450;
  wire [63:0] _result_T_1400 = _result_T_1398 + _result_T_451;
  wire [63:0] _result_T_1402 = _result_T_1400 + _result_T_452;
  wire [63:0] _result_T_1404 = _result_T_1402 + _result_T_453;
  wire [63:0] _result_T_1406 = _result_T_1404 + _result_T_454;
  wire [63:0] _result_T_1408 = _result_T_1406 + _result_T_455;
  wire [63:0] _result_T_1410 = _result_T_1408 + _result_T_456;
  wire [63:0] _result_T_1412 = _result_T_1410 + _result_T_457;
  wire [63:0] _result_T_1414 = _result_T_1412 + _result_T_458;
  wire [63:0] _result_T_1416 = _result_T_1414 + _result_T_459;
  wire [63:0] _result_T_1418 = _result_T_1416 + _result_T_460;
  wire [63:0] _result_T_1420 = _result_T_1418 + _result_T_461;
  wire [63:0] _result_T_1422 = _result_T_1420 + _result_T_462;
  wire [63:0] _result_T_1424 = _result_T_1422 + _result_T_463;
  wire [63:0] _result_T_1426 = _result_T_1424 + _result_T_464;
  wire [63:0] _result_T_1428 = _result_T_1426 + _result_T_465;
  wire [63:0] _result_T_1430 = _result_T_1428 + _result_T_466;
  wire [63:0] _result_T_1432 = _result_T_1430 + _result_T_467;
  wire [63:0] _result_T_1434 = _result_T_1432 + _result_T_468;
  wire [63:0] _result_T_1436 = _result_T_1434 + _result_T_469;
  wire [63:0] _result_T_1438 = _result_T_1436 + _result_T_470;
  wire [63:0] _result_T_1440 = _result_T_1438 + _result_T_471;
  wire [63:0] _result_T_1442 = _result_T_1440 + _result_T_472;
  wire [63:0] _result_T_1444 = _result_T_1442 + _result_T_473;
  wire [63:0] _result_T_1446 = _result_T_1444 + _result_T_474;
  wire [63:0] _result_T_1448 = _result_T_1446 + _result_T_475;
  wire [63:0] _result_T_1450 = _result_T_1448 + _result_T_476;
  wire [63:0] _result_T_1452 = _result_T_1450 + _result_T_477;
  wire [63:0] _result_T_1454 = _result_T_1452 + _result_T_478;
  wire [63:0] _result_T_1456 = _result_T_1454 + _result_T_479;
  wire [63:0] _result_T_1458 = _result_T_1456 + _result_T_480;
  wire [63:0] _result_T_1460 = _result_T_1458 + _result_T_481;
  wire [63:0] _result_T_1462 = _result_T_1460 + _result_T_482;
  wire [63:0] _result_T_1464 = _result_T_1462 + _result_T_483;
  wire [63:0] _result_T_1466 = _result_T_1464 + _result_T_484;
  wire [63:0] _result_T_1468 = _result_T_1466 + _result_T_485;
  wire [63:0] _result_T_1470 = _result_T_1468 + _result_T_486;
  wire [63:0] _result_T_1472 = _result_T_1470 + _result_T_487;
  wire [63:0] _result_T_1474 = _result_T_1472 + _result_T_488;
  wire [63:0] _result_T_1476 = _result_T_1474 + _result_T_489;
  wire [63:0] _result_T_1478 = _result_T_1476 + _result_T_490;
  wire [63:0] _result_T_1480 = _result_T_1478 + _result_T_491;
  wire [63:0] _result_T_1482 = _result_T_1480 + _result_T_492;
  wire [63:0] _result_T_1484 = _result_T_1482 + _result_T_493;
  wire [63:0] _result_T_1486 = _result_T_1484 + _result_T_494;
  wire [63:0] _result_T_1488 = _result_T_1486 + _result_T_495;
  wire [63:0] _result_T_1490 = _result_T_1488 + _result_T_496;
  wire [63:0] _result_T_1492 = _result_T_1490 + _result_T_497;
  wire [63:0] _result_T_1494 = _result_T_1492 + _result_T_498;
  wire [63:0] _result_T_1496 = _result_T_1494 + _result_T_499;
  wire [63:0] _result_T_1498 = _result_T_1496 + _result_T_500;
  wire [63:0] _GEN_1000 = insn[6:0] == 7'h3b ? _result_T_1498 : result;
  assign rd = result[31:0];
  always @(posedge clock) begin
    if (reset) begin
      coeffs_0 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h0 == rs2[8:0]) begin
          coeffs_0 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_1 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1 == rs2[8:0]) begin
          coeffs_1 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_2 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h2 == rs2[8:0]) begin
          coeffs_2 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_3 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h3 == rs2[8:0]) begin
          coeffs_3 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_4 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h4 == rs2[8:0]) begin
          coeffs_4 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_5 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h5 == rs2[8:0]) begin
          coeffs_5 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_6 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h6 == rs2[8:0]) begin
          coeffs_6 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_7 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h7 == rs2[8:0]) begin
          coeffs_7 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_8 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h8 == rs2[8:0]) begin
          coeffs_8 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_9 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h9 == rs2[8:0]) begin
          coeffs_9 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_10 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'ha == rs2[8:0]) begin
          coeffs_10 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_11 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hb == rs2[8:0]) begin
          coeffs_11 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_12 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hc == rs2[8:0]) begin
          coeffs_12 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_13 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hd == rs2[8:0]) begin
          coeffs_13 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_14 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'he == rs2[8:0]) begin
          coeffs_14 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_15 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hf == rs2[8:0]) begin
          coeffs_15 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_16 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h10 == rs2[8:0]) begin
          coeffs_16 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_17 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h11 == rs2[8:0]) begin
          coeffs_17 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_18 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h12 == rs2[8:0]) begin
          coeffs_18 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_19 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h13 == rs2[8:0]) begin
          coeffs_19 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_20 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h14 == rs2[8:0]) begin
          coeffs_20 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_21 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h15 == rs2[8:0]) begin
          coeffs_21 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_22 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h16 == rs2[8:0]) begin
          coeffs_22 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_23 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h17 == rs2[8:0]) begin
          coeffs_23 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_24 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h18 == rs2[8:0]) begin
          coeffs_24 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_25 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h19 == rs2[8:0]) begin
          coeffs_25 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_26 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1a == rs2[8:0]) begin
          coeffs_26 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_27 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1b == rs2[8:0]) begin
          coeffs_27 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_28 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1c == rs2[8:0]) begin
          coeffs_28 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_29 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1d == rs2[8:0]) begin
          coeffs_29 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_30 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1e == rs2[8:0]) begin
          coeffs_30 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_31 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1f == rs2[8:0]) begin
          coeffs_31 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_32 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h20 == rs2[8:0]) begin
          coeffs_32 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_33 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h21 == rs2[8:0]) begin
          coeffs_33 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_34 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h22 == rs2[8:0]) begin
          coeffs_34 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_35 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h23 == rs2[8:0]) begin
          coeffs_35 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_36 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h24 == rs2[8:0]) begin
          coeffs_36 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_37 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h25 == rs2[8:0]) begin
          coeffs_37 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_38 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h26 == rs2[8:0]) begin
          coeffs_38 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_39 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h27 == rs2[8:0]) begin
          coeffs_39 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_40 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h28 == rs2[8:0]) begin
          coeffs_40 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_41 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h29 == rs2[8:0]) begin
          coeffs_41 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_42 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h2a == rs2[8:0]) begin
          coeffs_42 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_43 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h2b == rs2[8:0]) begin
          coeffs_43 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_44 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h2c == rs2[8:0]) begin
          coeffs_44 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_45 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h2d == rs2[8:0]) begin
          coeffs_45 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_46 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h2e == rs2[8:0]) begin
          coeffs_46 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_47 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h2f == rs2[8:0]) begin
          coeffs_47 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_48 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h30 == rs2[8:0]) begin
          coeffs_48 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_49 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h31 == rs2[8:0]) begin
          coeffs_49 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_50 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h32 == rs2[8:0]) begin
          coeffs_50 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_51 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h33 == rs2[8:0]) begin
          coeffs_51 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_52 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h34 == rs2[8:0]) begin
          coeffs_52 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_53 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h35 == rs2[8:0]) begin
          coeffs_53 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_54 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h36 == rs2[8:0]) begin
          coeffs_54 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_55 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h37 == rs2[8:0]) begin
          coeffs_55 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_56 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h38 == rs2[8:0]) begin
          coeffs_56 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_57 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h39 == rs2[8:0]) begin
          coeffs_57 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_58 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h3a == rs2[8:0]) begin
          coeffs_58 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_59 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h3b == rs2[8:0]) begin
          coeffs_59 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_60 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h3c == rs2[8:0]) begin
          coeffs_60 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_61 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h3d == rs2[8:0]) begin
          coeffs_61 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_62 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h3e == rs2[8:0]) begin
          coeffs_62 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_63 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h3f == rs2[8:0]) begin
          coeffs_63 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_64 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h40 == rs2[8:0]) begin
          coeffs_64 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_65 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h41 == rs2[8:0]) begin
          coeffs_65 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_66 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h42 == rs2[8:0]) begin
          coeffs_66 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_67 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h43 == rs2[8:0]) begin
          coeffs_67 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_68 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h44 == rs2[8:0]) begin
          coeffs_68 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_69 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h45 == rs2[8:0]) begin
          coeffs_69 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_70 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h46 == rs2[8:0]) begin
          coeffs_70 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_71 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h47 == rs2[8:0]) begin
          coeffs_71 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_72 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h48 == rs2[8:0]) begin
          coeffs_72 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_73 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h49 == rs2[8:0]) begin
          coeffs_73 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_74 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h4a == rs2[8:0]) begin
          coeffs_74 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_75 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h4b == rs2[8:0]) begin
          coeffs_75 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_76 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h4c == rs2[8:0]) begin
          coeffs_76 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_77 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h4d == rs2[8:0]) begin
          coeffs_77 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_78 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h4e == rs2[8:0]) begin
          coeffs_78 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_79 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h4f == rs2[8:0]) begin
          coeffs_79 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_80 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h50 == rs2[8:0]) begin
          coeffs_80 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_81 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h51 == rs2[8:0]) begin
          coeffs_81 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_82 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h52 == rs2[8:0]) begin
          coeffs_82 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_83 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h53 == rs2[8:0]) begin
          coeffs_83 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_84 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h54 == rs2[8:0]) begin
          coeffs_84 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_85 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h55 == rs2[8:0]) begin
          coeffs_85 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_86 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h56 == rs2[8:0]) begin
          coeffs_86 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_87 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h57 == rs2[8:0]) begin
          coeffs_87 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_88 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h58 == rs2[8:0]) begin
          coeffs_88 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_89 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h59 == rs2[8:0]) begin
          coeffs_89 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_90 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h5a == rs2[8:0]) begin
          coeffs_90 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_91 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h5b == rs2[8:0]) begin
          coeffs_91 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_92 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h5c == rs2[8:0]) begin
          coeffs_92 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_93 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h5d == rs2[8:0]) begin
          coeffs_93 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_94 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h5e == rs2[8:0]) begin
          coeffs_94 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_95 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h5f == rs2[8:0]) begin
          coeffs_95 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_96 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h60 == rs2[8:0]) begin
          coeffs_96 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_97 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h61 == rs2[8:0]) begin
          coeffs_97 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_98 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h62 == rs2[8:0]) begin
          coeffs_98 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_99 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h63 == rs2[8:0]) begin
          coeffs_99 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_100 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h64 == rs2[8:0]) begin
          coeffs_100 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_101 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h65 == rs2[8:0]) begin
          coeffs_101 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_102 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h66 == rs2[8:0]) begin
          coeffs_102 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_103 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h67 == rs2[8:0]) begin
          coeffs_103 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_104 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h68 == rs2[8:0]) begin
          coeffs_104 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_105 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h69 == rs2[8:0]) begin
          coeffs_105 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_106 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h6a == rs2[8:0]) begin
          coeffs_106 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_107 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h6b == rs2[8:0]) begin
          coeffs_107 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_108 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h6c == rs2[8:0]) begin
          coeffs_108 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_109 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h6d == rs2[8:0]) begin
          coeffs_109 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_110 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h6e == rs2[8:0]) begin
          coeffs_110 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_111 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h6f == rs2[8:0]) begin
          coeffs_111 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_112 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h70 == rs2[8:0]) begin
          coeffs_112 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_113 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h71 == rs2[8:0]) begin
          coeffs_113 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_114 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h72 == rs2[8:0]) begin
          coeffs_114 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_115 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h73 == rs2[8:0]) begin
          coeffs_115 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_116 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h74 == rs2[8:0]) begin
          coeffs_116 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_117 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h75 == rs2[8:0]) begin
          coeffs_117 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_118 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h76 == rs2[8:0]) begin
          coeffs_118 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_119 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h77 == rs2[8:0]) begin
          coeffs_119 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_120 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h78 == rs2[8:0]) begin
          coeffs_120 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_121 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h79 == rs2[8:0]) begin
          coeffs_121 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_122 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h7a == rs2[8:0]) begin
          coeffs_122 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_123 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h7b == rs2[8:0]) begin
          coeffs_123 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_124 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h7c == rs2[8:0]) begin
          coeffs_124 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_125 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h7d == rs2[8:0]) begin
          coeffs_125 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_126 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h7e == rs2[8:0]) begin
          coeffs_126 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_127 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h7f == rs2[8:0]) begin
          coeffs_127 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_128 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h80 == rs2[8:0]) begin
          coeffs_128 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_129 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h81 == rs2[8:0]) begin
          coeffs_129 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_130 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h82 == rs2[8:0]) begin
          coeffs_130 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_131 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h83 == rs2[8:0]) begin
          coeffs_131 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_132 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h84 == rs2[8:0]) begin
          coeffs_132 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_133 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h85 == rs2[8:0]) begin
          coeffs_133 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_134 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h86 == rs2[8:0]) begin
          coeffs_134 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_135 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h87 == rs2[8:0]) begin
          coeffs_135 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_136 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h88 == rs2[8:0]) begin
          coeffs_136 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_137 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h89 == rs2[8:0]) begin
          coeffs_137 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_138 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h8a == rs2[8:0]) begin
          coeffs_138 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_139 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h8b == rs2[8:0]) begin
          coeffs_139 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_140 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h8c == rs2[8:0]) begin
          coeffs_140 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_141 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h8d == rs2[8:0]) begin
          coeffs_141 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_142 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h8e == rs2[8:0]) begin
          coeffs_142 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_143 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h8f == rs2[8:0]) begin
          coeffs_143 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_144 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h90 == rs2[8:0]) begin
          coeffs_144 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_145 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h91 == rs2[8:0]) begin
          coeffs_145 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_146 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h92 == rs2[8:0]) begin
          coeffs_146 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_147 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h93 == rs2[8:0]) begin
          coeffs_147 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_148 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h94 == rs2[8:0]) begin
          coeffs_148 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_149 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h95 == rs2[8:0]) begin
          coeffs_149 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_150 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h96 == rs2[8:0]) begin
          coeffs_150 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_151 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h97 == rs2[8:0]) begin
          coeffs_151 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_152 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h98 == rs2[8:0]) begin
          coeffs_152 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_153 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h99 == rs2[8:0]) begin
          coeffs_153 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_154 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h9a == rs2[8:0]) begin
          coeffs_154 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_155 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h9b == rs2[8:0]) begin
          coeffs_155 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_156 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h9c == rs2[8:0]) begin
          coeffs_156 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_157 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h9d == rs2[8:0]) begin
          coeffs_157 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_158 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h9e == rs2[8:0]) begin
          coeffs_158 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_159 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h9f == rs2[8:0]) begin
          coeffs_159 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_160 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'ha0 == rs2[8:0]) begin
          coeffs_160 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_161 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'ha1 == rs2[8:0]) begin
          coeffs_161 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_162 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'ha2 == rs2[8:0]) begin
          coeffs_162 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_163 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'ha3 == rs2[8:0]) begin
          coeffs_163 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_164 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'ha4 == rs2[8:0]) begin
          coeffs_164 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_165 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'ha5 == rs2[8:0]) begin
          coeffs_165 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_166 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'ha6 == rs2[8:0]) begin
          coeffs_166 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_167 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'ha7 == rs2[8:0]) begin
          coeffs_167 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_168 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'ha8 == rs2[8:0]) begin
          coeffs_168 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_169 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'ha9 == rs2[8:0]) begin
          coeffs_169 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_170 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'haa == rs2[8:0]) begin
          coeffs_170 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_171 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hab == rs2[8:0]) begin
          coeffs_171 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_172 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hac == rs2[8:0]) begin
          coeffs_172 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_173 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'had == rs2[8:0]) begin
          coeffs_173 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_174 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hae == rs2[8:0]) begin
          coeffs_174 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_175 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'haf == rs2[8:0]) begin
          coeffs_175 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_176 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hb0 == rs2[8:0]) begin
          coeffs_176 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_177 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hb1 == rs2[8:0]) begin
          coeffs_177 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_178 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hb2 == rs2[8:0]) begin
          coeffs_178 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_179 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hb3 == rs2[8:0]) begin
          coeffs_179 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_180 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hb4 == rs2[8:0]) begin
          coeffs_180 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_181 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hb5 == rs2[8:0]) begin
          coeffs_181 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_182 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hb6 == rs2[8:0]) begin
          coeffs_182 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_183 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hb7 == rs2[8:0]) begin
          coeffs_183 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_184 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hb8 == rs2[8:0]) begin
          coeffs_184 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_185 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hb9 == rs2[8:0]) begin
          coeffs_185 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_186 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hba == rs2[8:0]) begin
          coeffs_186 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_187 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hbb == rs2[8:0]) begin
          coeffs_187 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_188 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hbc == rs2[8:0]) begin
          coeffs_188 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_189 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hbd == rs2[8:0]) begin
          coeffs_189 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_190 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hbe == rs2[8:0]) begin
          coeffs_190 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_191 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hbf == rs2[8:0]) begin
          coeffs_191 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_192 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hc0 == rs2[8:0]) begin
          coeffs_192 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_193 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hc1 == rs2[8:0]) begin
          coeffs_193 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_194 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hc2 == rs2[8:0]) begin
          coeffs_194 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_195 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hc3 == rs2[8:0]) begin
          coeffs_195 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_196 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hc4 == rs2[8:0]) begin
          coeffs_196 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_197 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hc5 == rs2[8:0]) begin
          coeffs_197 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_198 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hc6 == rs2[8:0]) begin
          coeffs_198 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_199 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hc7 == rs2[8:0]) begin
          coeffs_199 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_200 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hc8 == rs2[8:0]) begin
          coeffs_200 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_201 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hc9 == rs2[8:0]) begin
          coeffs_201 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_202 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hca == rs2[8:0]) begin
          coeffs_202 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_203 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hcb == rs2[8:0]) begin
          coeffs_203 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_204 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hcc == rs2[8:0]) begin
          coeffs_204 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_205 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hcd == rs2[8:0]) begin
          coeffs_205 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_206 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hce == rs2[8:0]) begin
          coeffs_206 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_207 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hcf == rs2[8:0]) begin
          coeffs_207 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_208 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hd0 == rs2[8:0]) begin
          coeffs_208 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_209 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hd1 == rs2[8:0]) begin
          coeffs_209 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_210 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hd2 == rs2[8:0]) begin
          coeffs_210 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_211 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hd3 == rs2[8:0]) begin
          coeffs_211 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_212 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hd4 == rs2[8:0]) begin
          coeffs_212 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_213 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hd5 == rs2[8:0]) begin
          coeffs_213 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_214 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hd6 == rs2[8:0]) begin
          coeffs_214 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_215 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hd7 == rs2[8:0]) begin
          coeffs_215 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_216 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hd8 == rs2[8:0]) begin
          coeffs_216 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_217 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hd9 == rs2[8:0]) begin
          coeffs_217 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_218 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hda == rs2[8:0]) begin
          coeffs_218 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_219 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hdb == rs2[8:0]) begin
          coeffs_219 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_220 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hdc == rs2[8:0]) begin
          coeffs_220 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_221 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hdd == rs2[8:0]) begin
          coeffs_221 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_222 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hde == rs2[8:0]) begin
          coeffs_222 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_223 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hdf == rs2[8:0]) begin
          coeffs_223 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_224 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'he0 == rs2[8:0]) begin
          coeffs_224 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_225 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'he1 == rs2[8:0]) begin
          coeffs_225 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_226 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'he2 == rs2[8:0]) begin
          coeffs_226 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_227 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'he3 == rs2[8:0]) begin
          coeffs_227 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_228 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'he4 == rs2[8:0]) begin
          coeffs_228 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_229 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'he5 == rs2[8:0]) begin
          coeffs_229 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_230 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'he6 == rs2[8:0]) begin
          coeffs_230 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_231 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'he7 == rs2[8:0]) begin
          coeffs_231 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_232 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'he8 == rs2[8:0]) begin
          coeffs_232 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_233 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'he9 == rs2[8:0]) begin
          coeffs_233 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_234 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hea == rs2[8:0]) begin
          coeffs_234 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_235 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'heb == rs2[8:0]) begin
          coeffs_235 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_236 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hec == rs2[8:0]) begin
          coeffs_236 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_237 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hed == rs2[8:0]) begin
          coeffs_237 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_238 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hee == rs2[8:0]) begin
          coeffs_238 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_239 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hef == rs2[8:0]) begin
          coeffs_239 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_240 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hf0 == rs2[8:0]) begin
          coeffs_240 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_241 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hf1 == rs2[8:0]) begin
          coeffs_241 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_242 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hf2 == rs2[8:0]) begin
          coeffs_242 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_243 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hf3 == rs2[8:0]) begin
          coeffs_243 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_244 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hf4 == rs2[8:0]) begin
          coeffs_244 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_245 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hf5 == rs2[8:0]) begin
          coeffs_245 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_246 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hf6 == rs2[8:0]) begin
          coeffs_246 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_247 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hf7 == rs2[8:0]) begin
          coeffs_247 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_248 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hf8 == rs2[8:0]) begin
          coeffs_248 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_249 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hf9 == rs2[8:0]) begin
          coeffs_249 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_250 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hfa == rs2[8:0]) begin
          coeffs_250 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_251 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hfb == rs2[8:0]) begin
          coeffs_251 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_252 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hfc == rs2[8:0]) begin
          coeffs_252 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_253 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hfd == rs2[8:0]) begin
          coeffs_253 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_254 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hfe == rs2[8:0]) begin
          coeffs_254 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_255 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'hff == rs2[8:0]) begin
          coeffs_255 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_256 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h100 == rs2[8:0]) begin
          coeffs_256 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_257 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h101 == rs2[8:0]) begin
          coeffs_257 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_258 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h102 == rs2[8:0]) begin
          coeffs_258 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_259 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h103 == rs2[8:0]) begin
          coeffs_259 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_260 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h104 == rs2[8:0]) begin
          coeffs_260 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_261 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h105 == rs2[8:0]) begin
          coeffs_261 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_262 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h106 == rs2[8:0]) begin
          coeffs_262 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_263 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h107 == rs2[8:0]) begin
          coeffs_263 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_264 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h108 == rs2[8:0]) begin
          coeffs_264 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_265 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h109 == rs2[8:0]) begin
          coeffs_265 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_266 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h10a == rs2[8:0]) begin
          coeffs_266 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_267 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h10b == rs2[8:0]) begin
          coeffs_267 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_268 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h10c == rs2[8:0]) begin
          coeffs_268 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_269 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h10d == rs2[8:0]) begin
          coeffs_269 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_270 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h10e == rs2[8:0]) begin
          coeffs_270 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_271 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h10f == rs2[8:0]) begin
          coeffs_271 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_272 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h110 == rs2[8:0]) begin
          coeffs_272 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_273 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h111 == rs2[8:0]) begin
          coeffs_273 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_274 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h112 == rs2[8:0]) begin
          coeffs_274 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_275 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h113 == rs2[8:0]) begin
          coeffs_275 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_276 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h114 == rs2[8:0]) begin
          coeffs_276 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_277 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h115 == rs2[8:0]) begin
          coeffs_277 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_278 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h116 == rs2[8:0]) begin
          coeffs_278 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_279 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h117 == rs2[8:0]) begin
          coeffs_279 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_280 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h118 == rs2[8:0]) begin
          coeffs_280 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_281 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h119 == rs2[8:0]) begin
          coeffs_281 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_282 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h11a == rs2[8:0]) begin
          coeffs_282 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_283 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h11b == rs2[8:0]) begin
          coeffs_283 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_284 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h11c == rs2[8:0]) begin
          coeffs_284 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_285 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h11d == rs2[8:0]) begin
          coeffs_285 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_286 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h11e == rs2[8:0]) begin
          coeffs_286 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_287 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h11f == rs2[8:0]) begin
          coeffs_287 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_288 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h120 == rs2[8:0]) begin
          coeffs_288 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_289 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h121 == rs2[8:0]) begin
          coeffs_289 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_290 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h122 == rs2[8:0]) begin
          coeffs_290 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_291 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h123 == rs2[8:0]) begin
          coeffs_291 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_292 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h124 == rs2[8:0]) begin
          coeffs_292 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_293 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h125 == rs2[8:0]) begin
          coeffs_293 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_294 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h126 == rs2[8:0]) begin
          coeffs_294 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_295 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h127 == rs2[8:0]) begin
          coeffs_295 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_296 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h128 == rs2[8:0]) begin
          coeffs_296 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_297 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h129 == rs2[8:0]) begin
          coeffs_297 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_298 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h12a == rs2[8:0]) begin
          coeffs_298 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_299 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h12b == rs2[8:0]) begin
          coeffs_299 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_300 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h12c == rs2[8:0]) begin
          coeffs_300 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_301 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h12d == rs2[8:0]) begin
          coeffs_301 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_302 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h12e == rs2[8:0]) begin
          coeffs_302 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_303 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h12f == rs2[8:0]) begin
          coeffs_303 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_304 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h130 == rs2[8:0]) begin
          coeffs_304 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_305 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h131 == rs2[8:0]) begin
          coeffs_305 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_306 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h132 == rs2[8:0]) begin
          coeffs_306 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_307 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h133 == rs2[8:0]) begin
          coeffs_307 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_308 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h134 == rs2[8:0]) begin
          coeffs_308 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_309 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h135 == rs2[8:0]) begin
          coeffs_309 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_310 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h136 == rs2[8:0]) begin
          coeffs_310 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_311 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h137 == rs2[8:0]) begin
          coeffs_311 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_312 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h138 == rs2[8:0]) begin
          coeffs_312 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_313 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h139 == rs2[8:0]) begin
          coeffs_313 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_314 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h13a == rs2[8:0]) begin
          coeffs_314 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_315 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h13b == rs2[8:0]) begin
          coeffs_315 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_316 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h13c == rs2[8:0]) begin
          coeffs_316 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_317 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h13d == rs2[8:0]) begin
          coeffs_317 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_318 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h13e == rs2[8:0]) begin
          coeffs_318 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_319 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h13f == rs2[8:0]) begin
          coeffs_319 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_320 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h140 == rs2[8:0]) begin
          coeffs_320 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_321 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h141 == rs2[8:0]) begin
          coeffs_321 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_322 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h142 == rs2[8:0]) begin
          coeffs_322 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_323 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h143 == rs2[8:0]) begin
          coeffs_323 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_324 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h144 == rs2[8:0]) begin
          coeffs_324 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_325 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h145 == rs2[8:0]) begin
          coeffs_325 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_326 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h146 == rs2[8:0]) begin
          coeffs_326 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_327 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h147 == rs2[8:0]) begin
          coeffs_327 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_328 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h148 == rs2[8:0]) begin
          coeffs_328 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_329 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h149 == rs2[8:0]) begin
          coeffs_329 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_330 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h14a == rs2[8:0]) begin
          coeffs_330 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_331 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h14b == rs2[8:0]) begin
          coeffs_331 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_332 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h14c == rs2[8:0]) begin
          coeffs_332 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_333 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h14d == rs2[8:0]) begin
          coeffs_333 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_334 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h14e == rs2[8:0]) begin
          coeffs_334 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_335 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h14f == rs2[8:0]) begin
          coeffs_335 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_336 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h150 == rs2[8:0]) begin
          coeffs_336 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_337 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h151 == rs2[8:0]) begin
          coeffs_337 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_338 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h152 == rs2[8:0]) begin
          coeffs_338 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_339 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h153 == rs2[8:0]) begin
          coeffs_339 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_340 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h154 == rs2[8:0]) begin
          coeffs_340 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_341 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h155 == rs2[8:0]) begin
          coeffs_341 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_342 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h156 == rs2[8:0]) begin
          coeffs_342 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_343 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h157 == rs2[8:0]) begin
          coeffs_343 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_344 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h158 == rs2[8:0]) begin
          coeffs_344 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_345 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h159 == rs2[8:0]) begin
          coeffs_345 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_346 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h15a == rs2[8:0]) begin
          coeffs_346 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_347 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h15b == rs2[8:0]) begin
          coeffs_347 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_348 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h15c == rs2[8:0]) begin
          coeffs_348 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_349 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h15d == rs2[8:0]) begin
          coeffs_349 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_350 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h15e == rs2[8:0]) begin
          coeffs_350 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_351 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h15f == rs2[8:0]) begin
          coeffs_351 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_352 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h160 == rs2[8:0]) begin
          coeffs_352 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_353 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h161 == rs2[8:0]) begin
          coeffs_353 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_354 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h162 == rs2[8:0]) begin
          coeffs_354 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_355 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h163 == rs2[8:0]) begin
          coeffs_355 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_356 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h164 == rs2[8:0]) begin
          coeffs_356 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_357 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h165 == rs2[8:0]) begin
          coeffs_357 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_358 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h166 == rs2[8:0]) begin
          coeffs_358 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_359 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h167 == rs2[8:0]) begin
          coeffs_359 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_360 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h168 == rs2[8:0]) begin
          coeffs_360 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_361 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h169 == rs2[8:0]) begin
          coeffs_361 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_362 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h16a == rs2[8:0]) begin
          coeffs_362 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_363 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h16b == rs2[8:0]) begin
          coeffs_363 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_364 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h16c == rs2[8:0]) begin
          coeffs_364 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_365 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h16d == rs2[8:0]) begin
          coeffs_365 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_366 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h16e == rs2[8:0]) begin
          coeffs_366 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_367 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h16f == rs2[8:0]) begin
          coeffs_367 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_368 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h170 == rs2[8:0]) begin
          coeffs_368 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_369 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h171 == rs2[8:0]) begin
          coeffs_369 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_370 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h172 == rs2[8:0]) begin
          coeffs_370 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_371 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h173 == rs2[8:0]) begin
          coeffs_371 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_372 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h174 == rs2[8:0]) begin
          coeffs_372 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_373 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h175 == rs2[8:0]) begin
          coeffs_373 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_374 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h176 == rs2[8:0]) begin
          coeffs_374 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_375 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h177 == rs2[8:0]) begin
          coeffs_375 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_376 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h178 == rs2[8:0]) begin
          coeffs_376 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_377 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h179 == rs2[8:0]) begin
          coeffs_377 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_378 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h17a == rs2[8:0]) begin
          coeffs_378 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_379 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h17b == rs2[8:0]) begin
          coeffs_379 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_380 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h17c == rs2[8:0]) begin
          coeffs_380 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_381 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h17d == rs2[8:0]) begin
          coeffs_381 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_382 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h17e == rs2[8:0]) begin
          coeffs_382 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_383 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h17f == rs2[8:0]) begin
          coeffs_383 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_384 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h180 == rs2[8:0]) begin
          coeffs_384 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_385 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h181 == rs2[8:0]) begin
          coeffs_385 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_386 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h182 == rs2[8:0]) begin
          coeffs_386 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_387 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h183 == rs2[8:0]) begin
          coeffs_387 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_388 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h184 == rs2[8:0]) begin
          coeffs_388 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_389 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h185 == rs2[8:0]) begin
          coeffs_389 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_390 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h186 == rs2[8:0]) begin
          coeffs_390 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_391 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h187 == rs2[8:0]) begin
          coeffs_391 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_392 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h188 == rs2[8:0]) begin
          coeffs_392 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_393 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h189 == rs2[8:0]) begin
          coeffs_393 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_394 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h18a == rs2[8:0]) begin
          coeffs_394 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_395 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h18b == rs2[8:0]) begin
          coeffs_395 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_396 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h18c == rs2[8:0]) begin
          coeffs_396 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_397 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h18d == rs2[8:0]) begin
          coeffs_397 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_398 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h18e == rs2[8:0]) begin
          coeffs_398 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_399 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h18f == rs2[8:0]) begin
          coeffs_399 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_400 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h190 == rs2[8:0]) begin
          coeffs_400 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_401 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h191 == rs2[8:0]) begin
          coeffs_401 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_402 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h192 == rs2[8:0]) begin
          coeffs_402 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_403 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h193 == rs2[8:0]) begin
          coeffs_403 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_404 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h194 == rs2[8:0]) begin
          coeffs_404 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_405 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h195 == rs2[8:0]) begin
          coeffs_405 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_406 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h196 == rs2[8:0]) begin
          coeffs_406 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_407 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h197 == rs2[8:0]) begin
          coeffs_407 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_408 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h198 == rs2[8:0]) begin
          coeffs_408 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_409 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h199 == rs2[8:0]) begin
          coeffs_409 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_410 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h19a == rs2[8:0]) begin
          coeffs_410 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_411 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h19b == rs2[8:0]) begin
          coeffs_411 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_412 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h19c == rs2[8:0]) begin
          coeffs_412 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_413 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h19d == rs2[8:0]) begin
          coeffs_413 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_414 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h19e == rs2[8:0]) begin
          coeffs_414 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_415 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h19f == rs2[8:0]) begin
          coeffs_415 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_416 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1a0 == rs2[8:0]) begin
          coeffs_416 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_417 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1a1 == rs2[8:0]) begin
          coeffs_417 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_418 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1a2 == rs2[8:0]) begin
          coeffs_418 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_419 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1a3 == rs2[8:0]) begin
          coeffs_419 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_420 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1a4 == rs2[8:0]) begin
          coeffs_420 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_421 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1a5 == rs2[8:0]) begin
          coeffs_421 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_422 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1a6 == rs2[8:0]) begin
          coeffs_422 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_423 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1a7 == rs2[8:0]) begin
          coeffs_423 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_424 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1a8 == rs2[8:0]) begin
          coeffs_424 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_425 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1a9 == rs2[8:0]) begin
          coeffs_425 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_426 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1aa == rs2[8:0]) begin
          coeffs_426 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_427 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1ab == rs2[8:0]) begin
          coeffs_427 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_428 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1ac == rs2[8:0]) begin
          coeffs_428 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_429 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1ad == rs2[8:0]) begin
          coeffs_429 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_430 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1ae == rs2[8:0]) begin
          coeffs_430 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_431 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1af == rs2[8:0]) begin
          coeffs_431 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_432 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1b0 == rs2[8:0]) begin
          coeffs_432 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_433 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1b1 == rs2[8:0]) begin
          coeffs_433 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_434 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1b2 == rs2[8:0]) begin
          coeffs_434 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_435 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1b3 == rs2[8:0]) begin
          coeffs_435 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_436 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1b4 == rs2[8:0]) begin
          coeffs_436 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_437 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1b5 == rs2[8:0]) begin
          coeffs_437 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_438 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1b6 == rs2[8:0]) begin
          coeffs_438 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_439 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1b7 == rs2[8:0]) begin
          coeffs_439 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_440 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1b8 == rs2[8:0]) begin
          coeffs_440 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_441 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1b9 == rs2[8:0]) begin
          coeffs_441 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_442 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1ba == rs2[8:0]) begin
          coeffs_442 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_443 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1bb == rs2[8:0]) begin
          coeffs_443 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_444 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1bc == rs2[8:0]) begin
          coeffs_444 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_445 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1bd == rs2[8:0]) begin
          coeffs_445 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_446 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1be == rs2[8:0]) begin
          coeffs_446 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_447 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1bf == rs2[8:0]) begin
          coeffs_447 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_448 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1c0 == rs2[8:0]) begin
          coeffs_448 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_449 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1c1 == rs2[8:0]) begin
          coeffs_449 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_450 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1c2 == rs2[8:0]) begin
          coeffs_450 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_451 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1c3 == rs2[8:0]) begin
          coeffs_451 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_452 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1c4 == rs2[8:0]) begin
          coeffs_452 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_453 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1c5 == rs2[8:0]) begin
          coeffs_453 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_454 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1c6 == rs2[8:0]) begin
          coeffs_454 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_455 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1c7 == rs2[8:0]) begin
          coeffs_455 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_456 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1c8 == rs2[8:0]) begin
          coeffs_456 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_457 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1c9 == rs2[8:0]) begin
          coeffs_457 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_458 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1ca == rs2[8:0]) begin
          coeffs_458 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_459 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1cb == rs2[8:0]) begin
          coeffs_459 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_460 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1cc == rs2[8:0]) begin
          coeffs_460 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_461 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1cd == rs2[8:0]) begin
          coeffs_461 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_462 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1ce == rs2[8:0]) begin
          coeffs_462 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_463 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1cf == rs2[8:0]) begin
          coeffs_463 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_464 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1d0 == rs2[8:0]) begin
          coeffs_464 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_465 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1d1 == rs2[8:0]) begin
          coeffs_465 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_466 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1d2 == rs2[8:0]) begin
          coeffs_466 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_467 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1d3 == rs2[8:0]) begin
          coeffs_467 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_468 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1d4 == rs2[8:0]) begin
          coeffs_468 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_469 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1d5 == rs2[8:0]) begin
          coeffs_469 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_470 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1d6 == rs2[8:0]) begin
          coeffs_470 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_471 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1d7 == rs2[8:0]) begin
          coeffs_471 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_472 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1d8 == rs2[8:0]) begin
          coeffs_472 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_473 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1d9 == rs2[8:0]) begin
          coeffs_473 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_474 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1da == rs2[8:0]) begin
          coeffs_474 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_475 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1db == rs2[8:0]) begin
          coeffs_475 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_476 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1dc == rs2[8:0]) begin
          coeffs_476 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_477 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1dd == rs2[8:0]) begin
          coeffs_477 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_478 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1de == rs2[8:0]) begin
          coeffs_478 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_479 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1df == rs2[8:0]) begin
          coeffs_479 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_480 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1e0 == rs2[8:0]) begin
          coeffs_480 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_481 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1e1 == rs2[8:0]) begin
          coeffs_481 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_482 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1e2 == rs2[8:0]) begin
          coeffs_482 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_483 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1e3 == rs2[8:0]) begin
          coeffs_483 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_484 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1e4 == rs2[8:0]) begin
          coeffs_484 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_485 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1e5 == rs2[8:0]) begin
          coeffs_485 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_486 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1e6 == rs2[8:0]) begin
          coeffs_486 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_487 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1e7 == rs2[8:0]) begin
          coeffs_487 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_488 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1e8 == rs2[8:0]) begin
          coeffs_488 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_489 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1e9 == rs2[8:0]) begin
          coeffs_489 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_490 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1ea == rs2[8:0]) begin
          coeffs_490 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_491 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1eb == rs2[8:0]) begin
          coeffs_491 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_492 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1ec == rs2[8:0]) begin
          coeffs_492 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_493 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1ed == rs2[8:0]) begin
          coeffs_493 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_494 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1ee == rs2[8:0]) begin
          coeffs_494 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_495 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1ef == rs2[8:0]) begin
          coeffs_495 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_496 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1f0 == rs2[8:0]) begin
          coeffs_496 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_497 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1f1 == rs2[8:0]) begin
          coeffs_497 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_498 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1f2 == rs2[8:0]) begin
          coeffs_498 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_499 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (9'h1f3 == rs2[8:0]) begin
          coeffs_499 <= rs1;
        end
      end
    end
    if (reset) begin
      data_0 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_0 <= rs1;
        end
      end
    end
    if (reset) begin
      data_1 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_1 <= data_0;
        end
      end
    end
    if (reset) begin
      data_2 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_2 <= data_1;
        end
      end
    end
    if (reset) begin
      data_3 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_3 <= data_2;
        end
      end
    end
    if (reset) begin
      data_4 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_4 <= data_3;
        end
      end
    end
    if (reset) begin
      data_5 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_5 <= data_4;
        end
      end
    end
    if (reset) begin
      data_6 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_6 <= data_5;
        end
      end
    end
    if (reset) begin
      data_7 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_7 <= data_6;
        end
      end
    end
    if (reset) begin
      data_8 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_8 <= data_7;
        end
      end
    end
    if (reset) begin
      data_9 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_9 <= data_8;
        end
      end
    end
    if (reset) begin
      data_10 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_10 <= data_9;
        end
      end
    end
    if (reset) begin
      data_11 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_11 <= data_10;
        end
      end
    end
    if (reset) begin
      data_12 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_12 <= data_11;
        end
      end
    end
    if (reset) begin
      data_13 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_13 <= data_12;
        end
      end
    end
    if (reset) begin
      data_14 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_14 <= data_13;
        end
      end
    end
    if (reset) begin
      data_15 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_15 <= data_14;
        end
      end
    end
    if (reset) begin
      data_16 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_16 <= data_15;
        end
      end
    end
    if (reset) begin
      data_17 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_17 <= data_16;
        end
      end
    end
    if (reset) begin
      data_18 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_18 <= data_17;
        end
      end
    end
    if (reset) begin
      data_19 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_19 <= data_18;
        end
      end
    end
    if (reset) begin
      data_20 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_20 <= data_19;
        end
      end
    end
    if (reset) begin
      data_21 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_21 <= data_20;
        end
      end
    end
    if (reset) begin
      data_22 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_22 <= data_21;
        end
      end
    end
    if (reset) begin
      data_23 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_23 <= data_22;
        end
      end
    end
    if (reset) begin
      data_24 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_24 <= data_23;
        end
      end
    end
    if (reset) begin
      data_25 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_25 <= data_24;
        end
      end
    end
    if (reset) begin
      data_26 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_26 <= data_25;
        end
      end
    end
    if (reset) begin
      data_27 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_27 <= data_26;
        end
      end
    end
    if (reset) begin
      data_28 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_28 <= data_27;
        end
      end
    end
    if (reset) begin
      data_29 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_29 <= data_28;
        end
      end
    end
    if (reset) begin
      data_30 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_30 <= data_29;
        end
      end
    end
    if (reset) begin
      data_31 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_31 <= data_30;
        end
      end
    end
    if (reset) begin
      data_32 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_32 <= data_31;
        end
      end
    end
    if (reset) begin
      data_33 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_33 <= data_32;
        end
      end
    end
    if (reset) begin
      data_34 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_34 <= data_33;
        end
      end
    end
    if (reset) begin
      data_35 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_35 <= data_34;
        end
      end
    end
    if (reset) begin
      data_36 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_36 <= data_35;
        end
      end
    end
    if (reset) begin
      data_37 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_37 <= data_36;
        end
      end
    end
    if (reset) begin
      data_38 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_38 <= data_37;
        end
      end
    end
    if (reset) begin
      data_39 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_39 <= data_38;
        end
      end
    end
    if (reset) begin
      data_40 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_40 <= data_39;
        end
      end
    end
    if (reset) begin
      data_41 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_41 <= data_40;
        end
      end
    end
    if (reset) begin
      data_42 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_42 <= data_41;
        end
      end
    end
    if (reset) begin
      data_43 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_43 <= data_42;
        end
      end
    end
    if (reset) begin
      data_44 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_44 <= data_43;
        end
      end
    end
    if (reset) begin
      data_45 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_45 <= data_44;
        end
      end
    end
    if (reset) begin
      data_46 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_46 <= data_45;
        end
      end
    end
    if (reset) begin
      data_47 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_47 <= data_46;
        end
      end
    end
    if (reset) begin
      data_48 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_48 <= data_47;
        end
      end
    end
    if (reset) begin
      data_49 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_49 <= data_48;
        end
      end
    end
    if (reset) begin
      data_50 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_50 <= data_49;
        end
      end
    end
    if (reset) begin
      data_51 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_51 <= data_50;
        end
      end
    end
    if (reset) begin
      data_52 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_52 <= data_51;
        end
      end
    end
    if (reset) begin
      data_53 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_53 <= data_52;
        end
      end
    end
    if (reset) begin
      data_54 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_54 <= data_53;
        end
      end
    end
    if (reset) begin
      data_55 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_55 <= data_54;
        end
      end
    end
    if (reset) begin
      data_56 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_56 <= data_55;
        end
      end
    end
    if (reset) begin
      data_57 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_57 <= data_56;
        end
      end
    end
    if (reset) begin
      data_58 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_58 <= data_57;
        end
      end
    end
    if (reset) begin
      data_59 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_59 <= data_58;
        end
      end
    end
    if (reset) begin
      data_60 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_60 <= data_59;
        end
      end
    end
    if (reset) begin
      data_61 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_61 <= data_60;
        end
      end
    end
    if (reset) begin
      data_62 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_62 <= data_61;
        end
      end
    end
    if (reset) begin
      data_63 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_63 <= data_62;
        end
      end
    end
    if (reset) begin
      data_64 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_64 <= data_63;
        end
      end
    end
    if (reset) begin
      data_65 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_65 <= data_64;
        end
      end
    end
    if (reset) begin
      data_66 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_66 <= data_65;
        end
      end
    end
    if (reset) begin
      data_67 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_67 <= data_66;
        end
      end
    end
    if (reset) begin
      data_68 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_68 <= data_67;
        end
      end
    end
    if (reset) begin
      data_69 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_69 <= data_68;
        end
      end
    end
    if (reset) begin
      data_70 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_70 <= data_69;
        end
      end
    end
    if (reset) begin
      data_71 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_71 <= data_70;
        end
      end
    end
    if (reset) begin
      data_72 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_72 <= data_71;
        end
      end
    end
    if (reset) begin
      data_73 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_73 <= data_72;
        end
      end
    end
    if (reset) begin
      data_74 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_74 <= data_73;
        end
      end
    end
    if (reset) begin
      data_75 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_75 <= data_74;
        end
      end
    end
    if (reset) begin
      data_76 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_76 <= data_75;
        end
      end
    end
    if (reset) begin
      data_77 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_77 <= data_76;
        end
      end
    end
    if (reset) begin
      data_78 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_78 <= data_77;
        end
      end
    end
    if (reset) begin
      data_79 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_79 <= data_78;
        end
      end
    end
    if (reset) begin
      data_80 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_80 <= data_79;
        end
      end
    end
    if (reset) begin
      data_81 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_81 <= data_80;
        end
      end
    end
    if (reset) begin
      data_82 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_82 <= data_81;
        end
      end
    end
    if (reset) begin
      data_83 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_83 <= data_82;
        end
      end
    end
    if (reset) begin
      data_84 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_84 <= data_83;
        end
      end
    end
    if (reset) begin
      data_85 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_85 <= data_84;
        end
      end
    end
    if (reset) begin
      data_86 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_86 <= data_85;
        end
      end
    end
    if (reset) begin
      data_87 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_87 <= data_86;
        end
      end
    end
    if (reset) begin
      data_88 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_88 <= data_87;
        end
      end
    end
    if (reset) begin
      data_89 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_89 <= data_88;
        end
      end
    end
    if (reset) begin
      data_90 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_90 <= data_89;
        end
      end
    end
    if (reset) begin
      data_91 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_91 <= data_90;
        end
      end
    end
    if (reset) begin
      data_92 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_92 <= data_91;
        end
      end
    end
    if (reset) begin
      data_93 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_93 <= data_92;
        end
      end
    end
    if (reset) begin
      data_94 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_94 <= data_93;
        end
      end
    end
    if (reset) begin
      data_95 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_95 <= data_94;
        end
      end
    end
    if (reset) begin
      data_96 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_96 <= data_95;
        end
      end
    end
    if (reset) begin
      data_97 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_97 <= data_96;
        end
      end
    end
    if (reset) begin
      data_98 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_98 <= data_97;
        end
      end
    end
    if (reset) begin
      data_99 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_99 <= data_98;
        end
      end
    end
    if (reset) begin
      data_100 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_100 <= data_99;
        end
      end
    end
    if (reset) begin
      data_101 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_101 <= data_100;
        end
      end
    end
    if (reset) begin
      data_102 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_102 <= data_101;
        end
      end
    end
    if (reset) begin
      data_103 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_103 <= data_102;
        end
      end
    end
    if (reset) begin
      data_104 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_104 <= data_103;
        end
      end
    end
    if (reset) begin
      data_105 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_105 <= data_104;
        end
      end
    end
    if (reset) begin
      data_106 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_106 <= data_105;
        end
      end
    end
    if (reset) begin
      data_107 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_107 <= data_106;
        end
      end
    end
    if (reset) begin
      data_108 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_108 <= data_107;
        end
      end
    end
    if (reset) begin
      data_109 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_109 <= data_108;
        end
      end
    end
    if (reset) begin
      data_110 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_110 <= data_109;
        end
      end
    end
    if (reset) begin
      data_111 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_111 <= data_110;
        end
      end
    end
    if (reset) begin
      data_112 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_112 <= data_111;
        end
      end
    end
    if (reset) begin
      data_113 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_113 <= data_112;
        end
      end
    end
    if (reset) begin
      data_114 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_114 <= data_113;
        end
      end
    end
    if (reset) begin
      data_115 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_115 <= data_114;
        end
      end
    end
    if (reset) begin
      data_116 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_116 <= data_115;
        end
      end
    end
    if (reset) begin
      data_117 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_117 <= data_116;
        end
      end
    end
    if (reset) begin
      data_118 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_118 <= data_117;
        end
      end
    end
    if (reset) begin
      data_119 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_119 <= data_118;
        end
      end
    end
    if (reset) begin
      data_120 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_120 <= data_119;
        end
      end
    end
    if (reset) begin
      data_121 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_121 <= data_120;
        end
      end
    end
    if (reset) begin
      data_122 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_122 <= data_121;
        end
      end
    end
    if (reset) begin
      data_123 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_123 <= data_122;
        end
      end
    end
    if (reset) begin
      data_124 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_124 <= data_123;
        end
      end
    end
    if (reset) begin
      data_125 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_125 <= data_124;
        end
      end
    end
    if (reset) begin
      data_126 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_126 <= data_125;
        end
      end
    end
    if (reset) begin
      data_127 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_127 <= data_126;
        end
      end
    end
    if (reset) begin
      data_128 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_128 <= data_127;
        end
      end
    end
    if (reset) begin
      data_129 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_129 <= data_128;
        end
      end
    end
    if (reset) begin
      data_130 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_130 <= data_129;
        end
      end
    end
    if (reset) begin
      data_131 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_131 <= data_130;
        end
      end
    end
    if (reset) begin
      data_132 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_132 <= data_131;
        end
      end
    end
    if (reset) begin
      data_133 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_133 <= data_132;
        end
      end
    end
    if (reset) begin
      data_134 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_134 <= data_133;
        end
      end
    end
    if (reset) begin
      data_135 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_135 <= data_134;
        end
      end
    end
    if (reset) begin
      data_136 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_136 <= data_135;
        end
      end
    end
    if (reset) begin
      data_137 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_137 <= data_136;
        end
      end
    end
    if (reset) begin
      data_138 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_138 <= data_137;
        end
      end
    end
    if (reset) begin
      data_139 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_139 <= data_138;
        end
      end
    end
    if (reset) begin
      data_140 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_140 <= data_139;
        end
      end
    end
    if (reset) begin
      data_141 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_141 <= data_140;
        end
      end
    end
    if (reset) begin
      data_142 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_142 <= data_141;
        end
      end
    end
    if (reset) begin
      data_143 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_143 <= data_142;
        end
      end
    end
    if (reset) begin
      data_144 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_144 <= data_143;
        end
      end
    end
    if (reset) begin
      data_145 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_145 <= data_144;
        end
      end
    end
    if (reset) begin
      data_146 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_146 <= data_145;
        end
      end
    end
    if (reset) begin
      data_147 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_147 <= data_146;
        end
      end
    end
    if (reset) begin
      data_148 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_148 <= data_147;
        end
      end
    end
    if (reset) begin
      data_149 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_149 <= data_148;
        end
      end
    end
    if (reset) begin
      data_150 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_150 <= data_149;
        end
      end
    end
    if (reset) begin
      data_151 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_151 <= data_150;
        end
      end
    end
    if (reset) begin
      data_152 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_152 <= data_151;
        end
      end
    end
    if (reset) begin
      data_153 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_153 <= data_152;
        end
      end
    end
    if (reset) begin
      data_154 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_154 <= data_153;
        end
      end
    end
    if (reset) begin
      data_155 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_155 <= data_154;
        end
      end
    end
    if (reset) begin
      data_156 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_156 <= data_155;
        end
      end
    end
    if (reset) begin
      data_157 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_157 <= data_156;
        end
      end
    end
    if (reset) begin
      data_158 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_158 <= data_157;
        end
      end
    end
    if (reset) begin
      data_159 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_159 <= data_158;
        end
      end
    end
    if (reset) begin
      data_160 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_160 <= data_159;
        end
      end
    end
    if (reset) begin
      data_161 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_161 <= data_160;
        end
      end
    end
    if (reset) begin
      data_162 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_162 <= data_161;
        end
      end
    end
    if (reset) begin
      data_163 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_163 <= data_162;
        end
      end
    end
    if (reset) begin
      data_164 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_164 <= data_163;
        end
      end
    end
    if (reset) begin
      data_165 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_165 <= data_164;
        end
      end
    end
    if (reset) begin
      data_166 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_166 <= data_165;
        end
      end
    end
    if (reset) begin
      data_167 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_167 <= data_166;
        end
      end
    end
    if (reset) begin
      data_168 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_168 <= data_167;
        end
      end
    end
    if (reset) begin
      data_169 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_169 <= data_168;
        end
      end
    end
    if (reset) begin
      data_170 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_170 <= data_169;
        end
      end
    end
    if (reset) begin
      data_171 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_171 <= data_170;
        end
      end
    end
    if (reset) begin
      data_172 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_172 <= data_171;
        end
      end
    end
    if (reset) begin
      data_173 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_173 <= data_172;
        end
      end
    end
    if (reset) begin
      data_174 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_174 <= data_173;
        end
      end
    end
    if (reset) begin
      data_175 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_175 <= data_174;
        end
      end
    end
    if (reset) begin
      data_176 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_176 <= data_175;
        end
      end
    end
    if (reset) begin
      data_177 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_177 <= data_176;
        end
      end
    end
    if (reset) begin
      data_178 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_178 <= data_177;
        end
      end
    end
    if (reset) begin
      data_179 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_179 <= data_178;
        end
      end
    end
    if (reset) begin
      data_180 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_180 <= data_179;
        end
      end
    end
    if (reset) begin
      data_181 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_181 <= data_180;
        end
      end
    end
    if (reset) begin
      data_182 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_182 <= data_181;
        end
      end
    end
    if (reset) begin
      data_183 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_183 <= data_182;
        end
      end
    end
    if (reset) begin
      data_184 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_184 <= data_183;
        end
      end
    end
    if (reset) begin
      data_185 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_185 <= data_184;
        end
      end
    end
    if (reset) begin
      data_186 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_186 <= data_185;
        end
      end
    end
    if (reset) begin
      data_187 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_187 <= data_186;
        end
      end
    end
    if (reset) begin
      data_188 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_188 <= data_187;
        end
      end
    end
    if (reset) begin
      data_189 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_189 <= data_188;
        end
      end
    end
    if (reset) begin
      data_190 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_190 <= data_189;
        end
      end
    end
    if (reset) begin
      data_191 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_191 <= data_190;
        end
      end
    end
    if (reset) begin
      data_192 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_192 <= data_191;
        end
      end
    end
    if (reset) begin
      data_193 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_193 <= data_192;
        end
      end
    end
    if (reset) begin
      data_194 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_194 <= data_193;
        end
      end
    end
    if (reset) begin
      data_195 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_195 <= data_194;
        end
      end
    end
    if (reset) begin
      data_196 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_196 <= data_195;
        end
      end
    end
    if (reset) begin
      data_197 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_197 <= data_196;
        end
      end
    end
    if (reset) begin
      data_198 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_198 <= data_197;
        end
      end
    end
    if (reset) begin
      data_199 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_199 <= data_198;
        end
      end
    end
    if (reset) begin
      data_200 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_200 <= data_199;
        end
      end
    end
    if (reset) begin
      data_201 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_201 <= data_200;
        end
      end
    end
    if (reset) begin
      data_202 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_202 <= data_201;
        end
      end
    end
    if (reset) begin
      data_203 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_203 <= data_202;
        end
      end
    end
    if (reset) begin
      data_204 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_204 <= data_203;
        end
      end
    end
    if (reset) begin
      data_205 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_205 <= data_204;
        end
      end
    end
    if (reset) begin
      data_206 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_206 <= data_205;
        end
      end
    end
    if (reset) begin
      data_207 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_207 <= data_206;
        end
      end
    end
    if (reset) begin
      data_208 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_208 <= data_207;
        end
      end
    end
    if (reset) begin
      data_209 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_209 <= data_208;
        end
      end
    end
    if (reset) begin
      data_210 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_210 <= data_209;
        end
      end
    end
    if (reset) begin
      data_211 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_211 <= data_210;
        end
      end
    end
    if (reset) begin
      data_212 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_212 <= data_211;
        end
      end
    end
    if (reset) begin
      data_213 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_213 <= data_212;
        end
      end
    end
    if (reset) begin
      data_214 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_214 <= data_213;
        end
      end
    end
    if (reset) begin
      data_215 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_215 <= data_214;
        end
      end
    end
    if (reset) begin
      data_216 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_216 <= data_215;
        end
      end
    end
    if (reset) begin
      data_217 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_217 <= data_216;
        end
      end
    end
    if (reset) begin
      data_218 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_218 <= data_217;
        end
      end
    end
    if (reset) begin
      data_219 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_219 <= data_218;
        end
      end
    end
    if (reset) begin
      data_220 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_220 <= data_219;
        end
      end
    end
    if (reset) begin
      data_221 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_221 <= data_220;
        end
      end
    end
    if (reset) begin
      data_222 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_222 <= data_221;
        end
      end
    end
    if (reset) begin
      data_223 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_223 <= data_222;
        end
      end
    end
    if (reset) begin
      data_224 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_224 <= data_223;
        end
      end
    end
    if (reset) begin
      data_225 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_225 <= data_224;
        end
      end
    end
    if (reset) begin
      data_226 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_226 <= data_225;
        end
      end
    end
    if (reset) begin
      data_227 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_227 <= data_226;
        end
      end
    end
    if (reset) begin
      data_228 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_228 <= data_227;
        end
      end
    end
    if (reset) begin
      data_229 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_229 <= data_228;
        end
      end
    end
    if (reset) begin
      data_230 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_230 <= data_229;
        end
      end
    end
    if (reset) begin
      data_231 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_231 <= data_230;
        end
      end
    end
    if (reset) begin
      data_232 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_232 <= data_231;
        end
      end
    end
    if (reset) begin
      data_233 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_233 <= data_232;
        end
      end
    end
    if (reset) begin
      data_234 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_234 <= data_233;
        end
      end
    end
    if (reset) begin
      data_235 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_235 <= data_234;
        end
      end
    end
    if (reset) begin
      data_236 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_236 <= data_235;
        end
      end
    end
    if (reset) begin
      data_237 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_237 <= data_236;
        end
      end
    end
    if (reset) begin
      data_238 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_238 <= data_237;
        end
      end
    end
    if (reset) begin
      data_239 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_239 <= data_238;
        end
      end
    end
    if (reset) begin
      data_240 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_240 <= data_239;
        end
      end
    end
    if (reset) begin
      data_241 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_241 <= data_240;
        end
      end
    end
    if (reset) begin
      data_242 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_242 <= data_241;
        end
      end
    end
    if (reset) begin
      data_243 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_243 <= data_242;
        end
      end
    end
    if (reset) begin
      data_244 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_244 <= data_243;
        end
      end
    end
    if (reset) begin
      data_245 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_245 <= data_244;
        end
      end
    end
    if (reset) begin
      data_246 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_246 <= data_245;
        end
      end
    end
    if (reset) begin
      data_247 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_247 <= data_246;
        end
      end
    end
    if (reset) begin
      data_248 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_248 <= data_247;
        end
      end
    end
    if (reset) begin
      data_249 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_249 <= data_248;
        end
      end
    end
    if (reset) begin
      data_250 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_250 <= data_249;
        end
      end
    end
    if (reset) begin
      data_251 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_251 <= data_250;
        end
      end
    end
    if (reset) begin
      data_252 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_252 <= data_251;
        end
      end
    end
    if (reset) begin
      data_253 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_253 <= data_252;
        end
      end
    end
    if (reset) begin
      data_254 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_254 <= data_253;
        end
      end
    end
    if (reset) begin
      data_255 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_255 <= data_254;
        end
      end
    end
    if (reset) begin
      data_256 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_256 <= data_255;
        end
      end
    end
    if (reset) begin
      data_257 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_257 <= data_256;
        end
      end
    end
    if (reset) begin
      data_258 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_258 <= data_257;
        end
      end
    end
    if (reset) begin
      data_259 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_259 <= data_258;
        end
      end
    end
    if (reset) begin
      data_260 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_260 <= data_259;
        end
      end
    end
    if (reset) begin
      data_261 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_261 <= data_260;
        end
      end
    end
    if (reset) begin
      data_262 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_262 <= data_261;
        end
      end
    end
    if (reset) begin
      data_263 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_263 <= data_262;
        end
      end
    end
    if (reset) begin
      data_264 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_264 <= data_263;
        end
      end
    end
    if (reset) begin
      data_265 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_265 <= data_264;
        end
      end
    end
    if (reset) begin
      data_266 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_266 <= data_265;
        end
      end
    end
    if (reset) begin
      data_267 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_267 <= data_266;
        end
      end
    end
    if (reset) begin
      data_268 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_268 <= data_267;
        end
      end
    end
    if (reset) begin
      data_269 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_269 <= data_268;
        end
      end
    end
    if (reset) begin
      data_270 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_270 <= data_269;
        end
      end
    end
    if (reset) begin
      data_271 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_271 <= data_270;
        end
      end
    end
    if (reset) begin
      data_272 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_272 <= data_271;
        end
      end
    end
    if (reset) begin
      data_273 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_273 <= data_272;
        end
      end
    end
    if (reset) begin
      data_274 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_274 <= data_273;
        end
      end
    end
    if (reset) begin
      data_275 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_275 <= data_274;
        end
      end
    end
    if (reset) begin
      data_276 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_276 <= data_275;
        end
      end
    end
    if (reset) begin
      data_277 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_277 <= data_276;
        end
      end
    end
    if (reset) begin
      data_278 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_278 <= data_277;
        end
      end
    end
    if (reset) begin
      data_279 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_279 <= data_278;
        end
      end
    end
    if (reset) begin
      data_280 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_280 <= data_279;
        end
      end
    end
    if (reset) begin
      data_281 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_281 <= data_280;
        end
      end
    end
    if (reset) begin
      data_282 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_282 <= data_281;
        end
      end
    end
    if (reset) begin
      data_283 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_283 <= data_282;
        end
      end
    end
    if (reset) begin
      data_284 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_284 <= data_283;
        end
      end
    end
    if (reset) begin
      data_285 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_285 <= data_284;
        end
      end
    end
    if (reset) begin
      data_286 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_286 <= data_285;
        end
      end
    end
    if (reset) begin
      data_287 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_287 <= data_286;
        end
      end
    end
    if (reset) begin
      data_288 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_288 <= data_287;
        end
      end
    end
    if (reset) begin
      data_289 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_289 <= data_288;
        end
      end
    end
    if (reset) begin
      data_290 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_290 <= data_289;
        end
      end
    end
    if (reset) begin
      data_291 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_291 <= data_290;
        end
      end
    end
    if (reset) begin
      data_292 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_292 <= data_291;
        end
      end
    end
    if (reset) begin
      data_293 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_293 <= data_292;
        end
      end
    end
    if (reset) begin
      data_294 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_294 <= data_293;
        end
      end
    end
    if (reset) begin
      data_295 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_295 <= data_294;
        end
      end
    end
    if (reset) begin
      data_296 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_296 <= data_295;
        end
      end
    end
    if (reset) begin
      data_297 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_297 <= data_296;
        end
      end
    end
    if (reset) begin
      data_298 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_298 <= data_297;
        end
      end
    end
    if (reset) begin
      data_299 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_299 <= data_298;
        end
      end
    end
    if (reset) begin
      data_300 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_300 <= data_299;
        end
      end
    end
    if (reset) begin
      data_301 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_301 <= data_300;
        end
      end
    end
    if (reset) begin
      data_302 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_302 <= data_301;
        end
      end
    end
    if (reset) begin
      data_303 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_303 <= data_302;
        end
      end
    end
    if (reset) begin
      data_304 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_304 <= data_303;
        end
      end
    end
    if (reset) begin
      data_305 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_305 <= data_304;
        end
      end
    end
    if (reset) begin
      data_306 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_306 <= data_305;
        end
      end
    end
    if (reset) begin
      data_307 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_307 <= data_306;
        end
      end
    end
    if (reset) begin
      data_308 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_308 <= data_307;
        end
      end
    end
    if (reset) begin
      data_309 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_309 <= data_308;
        end
      end
    end
    if (reset) begin
      data_310 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_310 <= data_309;
        end
      end
    end
    if (reset) begin
      data_311 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_311 <= data_310;
        end
      end
    end
    if (reset) begin
      data_312 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_312 <= data_311;
        end
      end
    end
    if (reset) begin
      data_313 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_313 <= data_312;
        end
      end
    end
    if (reset) begin
      data_314 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_314 <= data_313;
        end
      end
    end
    if (reset) begin
      data_315 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_315 <= data_314;
        end
      end
    end
    if (reset) begin
      data_316 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_316 <= data_315;
        end
      end
    end
    if (reset) begin
      data_317 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_317 <= data_316;
        end
      end
    end
    if (reset) begin
      data_318 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_318 <= data_317;
        end
      end
    end
    if (reset) begin
      data_319 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_319 <= data_318;
        end
      end
    end
    if (reset) begin
      data_320 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_320 <= data_319;
        end
      end
    end
    if (reset) begin
      data_321 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_321 <= data_320;
        end
      end
    end
    if (reset) begin
      data_322 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_322 <= data_321;
        end
      end
    end
    if (reset) begin
      data_323 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_323 <= data_322;
        end
      end
    end
    if (reset) begin
      data_324 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_324 <= data_323;
        end
      end
    end
    if (reset) begin
      data_325 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_325 <= data_324;
        end
      end
    end
    if (reset) begin
      data_326 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_326 <= data_325;
        end
      end
    end
    if (reset) begin
      data_327 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_327 <= data_326;
        end
      end
    end
    if (reset) begin
      data_328 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_328 <= data_327;
        end
      end
    end
    if (reset) begin
      data_329 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_329 <= data_328;
        end
      end
    end
    if (reset) begin
      data_330 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_330 <= data_329;
        end
      end
    end
    if (reset) begin
      data_331 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_331 <= data_330;
        end
      end
    end
    if (reset) begin
      data_332 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_332 <= data_331;
        end
      end
    end
    if (reset) begin
      data_333 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_333 <= data_332;
        end
      end
    end
    if (reset) begin
      data_334 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_334 <= data_333;
        end
      end
    end
    if (reset) begin
      data_335 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_335 <= data_334;
        end
      end
    end
    if (reset) begin
      data_336 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_336 <= data_335;
        end
      end
    end
    if (reset) begin
      data_337 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_337 <= data_336;
        end
      end
    end
    if (reset) begin
      data_338 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_338 <= data_337;
        end
      end
    end
    if (reset) begin
      data_339 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_339 <= data_338;
        end
      end
    end
    if (reset) begin
      data_340 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_340 <= data_339;
        end
      end
    end
    if (reset) begin
      data_341 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_341 <= data_340;
        end
      end
    end
    if (reset) begin
      data_342 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_342 <= data_341;
        end
      end
    end
    if (reset) begin
      data_343 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_343 <= data_342;
        end
      end
    end
    if (reset) begin
      data_344 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_344 <= data_343;
        end
      end
    end
    if (reset) begin
      data_345 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_345 <= data_344;
        end
      end
    end
    if (reset) begin
      data_346 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_346 <= data_345;
        end
      end
    end
    if (reset) begin
      data_347 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_347 <= data_346;
        end
      end
    end
    if (reset) begin
      data_348 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_348 <= data_347;
        end
      end
    end
    if (reset) begin
      data_349 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_349 <= data_348;
        end
      end
    end
    if (reset) begin
      data_350 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_350 <= data_349;
        end
      end
    end
    if (reset) begin
      data_351 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_351 <= data_350;
        end
      end
    end
    if (reset) begin
      data_352 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_352 <= data_351;
        end
      end
    end
    if (reset) begin
      data_353 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_353 <= data_352;
        end
      end
    end
    if (reset) begin
      data_354 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_354 <= data_353;
        end
      end
    end
    if (reset) begin
      data_355 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_355 <= data_354;
        end
      end
    end
    if (reset) begin
      data_356 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_356 <= data_355;
        end
      end
    end
    if (reset) begin
      data_357 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_357 <= data_356;
        end
      end
    end
    if (reset) begin
      data_358 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_358 <= data_357;
        end
      end
    end
    if (reset) begin
      data_359 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_359 <= data_358;
        end
      end
    end
    if (reset) begin
      data_360 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_360 <= data_359;
        end
      end
    end
    if (reset) begin
      data_361 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_361 <= data_360;
        end
      end
    end
    if (reset) begin
      data_362 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_362 <= data_361;
        end
      end
    end
    if (reset) begin
      data_363 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_363 <= data_362;
        end
      end
    end
    if (reset) begin
      data_364 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_364 <= data_363;
        end
      end
    end
    if (reset) begin
      data_365 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_365 <= data_364;
        end
      end
    end
    if (reset) begin
      data_366 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_366 <= data_365;
        end
      end
    end
    if (reset) begin
      data_367 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_367 <= data_366;
        end
      end
    end
    if (reset) begin
      data_368 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_368 <= data_367;
        end
      end
    end
    if (reset) begin
      data_369 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_369 <= data_368;
        end
      end
    end
    if (reset) begin
      data_370 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_370 <= data_369;
        end
      end
    end
    if (reset) begin
      data_371 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_371 <= data_370;
        end
      end
    end
    if (reset) begin
      data_372 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_372 <= data_371;
        end
      end
    end
    if (reset) begin
      data_373 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_373 <= data_372;
        end
      end
    end
    if (reset) begin
      data_374 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_374 <= data_373;
        end
      end
    end
    if (reset) begin
      data_375 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_375 <= data_374;
        end
      end
    end
    if (reset) begin
      data_376 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_376 <= data_375;
        end
      end
    end
    if (reset) begin
      data_377 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_377 <= data_376;
        end
      end
    end
    if (reset) begin
      data_378 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_378 <= data_377;
        end
      end
    end
    if (reset) begin
      data_379 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_379 <= data_378;
        end
      end
    end
    if (reset) begin
      data_380 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_380 <= data_379;
        end
      end
    end
    if (reset) begin
      data_381 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_381 <= data_380;
        end
      end
    end
    if (reset) begin
      data_382 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_382 <= data_381;
        end
      end
    end
    if (reset) begin
      data_383 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_383 <= data_382;
        end
      end
    end
    if (reset) begin
      data_384 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_384 <= data_383;
        end
      end
    end
    if (reset) begin
      data_385 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_385 <= data_384;
        end
      end
    end
    if (reset) begin
      data_386 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_386 <= data_385;
        end
      end
    end
    if (reset) begin
      data_387 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_387 <= data_386;
        end
      end
    end
    if (reset) begin
      data_388 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_388 <= data_387;
        end
      end
    end
    if (reset) begin
      data_389 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_389 <= data_388;
        end
      end
    end
    if (reset) begin
      data_390 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_390 <= data_389;
        end
      end
    end
    if (reset) begin
      data_391 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_391 <= data_390;
        end
      end
    end
    if (reset) begin
      data_392 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_392 <= data_391;
        end
      end
    end
    if (reset) begin
      data_393 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_393 <= data_392;
        end
      end
    end
    if (reset) begin
      data_394 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_394 <= data_393;
        end
      end
    end
    if (reset) begin
      data_395 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_395 <= data_394;
        end
      end
    end
    if (reset) begin
      data_396 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_396 <= data_395;
        end
      end
    end
    if (reset) begin
      data_397 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_397 <= data_396;
        end
      end
    end
    if (reset) begin
      data_398 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_398 <= data_397;
        end
      end
    end
    if (reset) begin
      data_399 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_399 <= data_398;
        end
      end
    end
    if (reset) begin
      data_400 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_400 <= data_399;
        end
      end
    end
    if (reset) begin
      data_401 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_401 <= data_400;
        end
      end
    end
    if (reset) begin
      data_402 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_402 <= data_401;
        end
      end
    end
    if (reset) begin
      data_403 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_403 <= data_402;
        end
      end
    end
    if (reset) begin
      data_404 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_404 <= data_403;
        end
      end
    end
    if (reset) begin
      data_405 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_405 <= data_404;
        end
      end
    end
    if (reset) begin
      data_406 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_406 <= data_405;
        end
      end
    end
    if (reset) begin
      data_407 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_407 <= data_406;
        end
      end
    end
    if (reset) begin
      data_408 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_408 <= data_407;
        end
      end
    end
    if (reset) begin
      data_409 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_409 <= data_408;
        end
      end
    end
    if (reset) begin
      data_410 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_410 <= data_409;
        end
      end
    end
    if (reset) begin
      data_411 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_411 <= data_410;
        end
      end
    end
    if (reset) begin
      data_412 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_412 <= data_411;
        end
      end
    end
    if (reset) begin
      data_413 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_413 <= data_412;
        end
      end
    end
    if (reset) begin
      data_414 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_414 <= data_413;
        end
      end
    end
    if (reset) begin
      data_415 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_415 <= data_414;
        end
      end
    end
    if (reset) begin
      data_416 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_416 <= data_415;
        end
      end
    end
    if (reset) begin
      data_417 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_417 <= data_416;
        end
      end
    end
    if (reset) begin
      data_418 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_418 <= data_417;
        end
      end
    end
    if (reset) begin
      data_419 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_419 <= data_418;
        end
      end
    end
    if (reset) begin
      data_420 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_420 <= data_419;
        end
      end
    end
    if (reset) begin
      data_421 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_421 <= data_420;
        end
      end
    end
    if (reset) begin
      data_422 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_422 <= data_421;
        end
      end
    end
    if (reset) begin
      data_423 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_423 <= data_422;
        end
      end
    end
    if (reset) begin
      data_424 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_424 <= data_423;
        end
      end
    end
    if (reset) begin
      data_425 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_425 <= data_424;
        end
      end
    end
    if (reset) begin
      data_426 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_426 <= data_425;
        end
      end
    end
    if (reset) begin
      data_427 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_427 <= data_426;
        end
      end
    end
    if (reset) begin
      data_428 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_428 <= data_427;
        end
      end
    end
    if (reset) begin
      data_429 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_429 <= data_428;
        end
      end
    end
    if (reset) begin
      data_430 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_430 <= data_429;
        end
      end
    end
    if (reset) begin
      data_431 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_431 <= data_430;
        end
      end
    end
    if (reset) begin
      data_432 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_432 <= data_431;
        end
      end
    end
    if (reset) begin
      data_433 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_433 <= data_432;
        end
      end
    end
    if (reset) begin
      data_434 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_434 <= data_433;
        end
      end
    end
    if (reset) begin
      data_435 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_435 <= data_434;
        end
      end
    end
    if (reset) begin
      data_436 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_436 <= data_435;
        end
      end
    end
    if (reset) begin
      data_437 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_437 <= data_436;
        end
      end
    end
    if (reset) begin
      data_438 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_438 <= data_437;
        end
      end
    end
    if (reset) begin
      data_439 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_439 <= data_438;
        end
      end
    end
    if (reset) begin
      data_440 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_440 <= data_439;
        end
      end
    end
    if (reset) begin
      data_441 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_441 <= data_440;
        end
      end
    end
    if (reset) begin
      data_442 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_442 <= data_441;
        end
      end
    end
    if (reset) begin
      data_443 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_443 <= data_442;
        end
      end
    end
    if (reset) begin
      data_444 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_444 <= data_443;
        end
      end
    end
    if (reset) begin
      data_445 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_445 <= data_444;
        end
      end
    end
    if (reset) begin
      data_446 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_446 <= data_445;
        end
      end
    end
    if (reset) begin
      data_447 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_447 <= data_446;
        end
      end
    end
    if (reset) begin
      data_448 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_448 <= data_447;
        end
      end
    end
    if (reset) begin
      data_449 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_449 <= data_448;
        end
      end
    end
    if (reset) begin
      data_450 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_450 <= data_449;
        end
      end
    end
    if (reset) begin
      data_451 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_451 <= data_450;
        end
      end
    end
    if (reset) begin
      data_452 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_452 <= data_451;
        end
      end
    end
    if (reset) begin
      data_453 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_453 <= data_452;
        end
      end
    end
    if (reset) begin
      data_454 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_454 <= data_453;
        end
      end
    end
    if (reset) begin
      data_455 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_455 <= data_454;
        end
      end
    end
    if (reset) begin
      data_456 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_456 <= data_455;
        end
      end
    end
    if (reset) begin
      data_457 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_457 <= data_456;
        end
      end
    end
    if (reset) begin
      data_458 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_458 <= data_457;
        end
      end
    end
    if (reset) begin
      data_459 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_459 <= data_458;
        end
      end
    end
    if (reset) begin
      data_460 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_460 <= data_459;
        end
      end
    end
    if (reset) begin
      data_461 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_461 <= data_460;
        end
      end
    end
    if (reset) begin
      data_462 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_462 <= data_461;
        end
      end
    end
    if (reset) begin
      data_463 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_463 <= data_462;
        end
      end
    end
    if (reset) begin
      data_464 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_464 <= data_463;
        end
      end
    end
    if (reset) begin
      data_465 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_465 <= data_464;
        end
      end
    end
    if (reset) begin
      data_466 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_466 <= data_465;
        end
      end
    end
    if (reset) begin
      data_467 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_467 <= data_466;
        end
      end
    end
    if (reset) begin
      data_468 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_468 <= data_467;
        end
      end
    end
    if (reset) begin
      data_469 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_469 <= data_468;
        end
      end
    end
    if (reset) begin
      data_470 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_470 <= data_469;
        end
      end
    end
    if (reset) begin
      data_471 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_471 <= data_470;
        end
      end
    end
    if (reset) begin
      data_472 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_472 <= data_471;
        end
      end
    end
    if (reset) begin
      data_473 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_473 <= data_472;
        end
      end
    end
    if (reset) begin
      data_474 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_474 <= data_473;
        end
      end
    end
    if (reset) begin
      data_475 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_475 <= data_474;
        end
      end
    end
    if (reset) begin
      data_476 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_476 <= data_475;
        end
      end
    end
    if (reset) begin
      data_477 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_477 <= data_476;
        end
      end
    end
    if (reset) begin
      data_478 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_478 <= data_477;
        end
      end
    end
    if (reset) begin
      data_479 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_479 <= data_478;
        end
      end
    end
    if (reset) begin
      data_480 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_480 <= data_479;
        end
      end
    end
    if (reset) begin
      data_481 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_481 <= data_480;
        end
      end
    end
    if (reset) begin
      data_482 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_482 <= data_481;
        end
      end
    end
    if (reset) begin
      data_483 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_483 <= data_482;
        end
      end
    end
    if (reset) begin
      data_484 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_484 <= data_483;
        end
      end
    end
    if (reset) begin
      data_485 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_485 <= data_484;
        end
      end
    end
    if (reset) begin
      data_486 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_486 <= data_485;
        end
      end
    end
    if (reset) begin
      data_487 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_487 <= data_486;
        end
      end
    end
    if (reset) begin
      data_488 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_488 <= data_487;
        end
      end
    end
    if (reset) begin
      data_489 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_489 <= data_488;
        end
      end
    end
    if (reset) begin
      data_490 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_490 <= data_489;
        end
      end
    end
    if (reset) begin
      data_491 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_491 <= data_490;
        end
      end
    end
    if (reset) begin
      data_492 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_492 <= data_491;
        end
      end
    end
    if (reset) begin
      data_493 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_493 <= data_492;
        end
      end
    end
    if (reset) begin
      data_494 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_494 <= data_493;
        end
      end
    end
    if (reset) begin
      data_495 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_495 <= data_494;
        end
      end
    end
    if (reset) begin
      data_496 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_496 <= data_495;
        end
      end
    end
    if (reset) begin
      data_497 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_497 <= data_496;
        end
      end
    end
    if (reset) begin
      data_498 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_498 <= data_497;
        end
      end
    end
    if (reset) begin
      data_499 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_499 <= data_498;
        end
      end
    end
    if (reset) begin
      result <= 64'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        result <= {{32'd0}, _GEN_999};
      end else if (insn[6:0] == 7'h2b) begin
        result <= {{32'd0}, data_0};
      end else begin
        result <= _GEN_1000;
      end
    end
  end
endmodule
