module SCIEPipelined #(parameter XLEN = 32)(
  input         clock,
  input         reset,
  input         valid,
  input  [31:0] insn,
  input  [31:0] rs1,
  input  [31:0] rs2,
  output [31:0] rd
);
  reg [31:0] coeffs_0;
  reg [31:0] coeffs_1;
  reg [31:0] coeffs_2;
  reg [31:0] coeffs_3;
  reg [31:0] coeffs_4;
  reg [31:0] coeffs_5;
  reg [31:0] coeffs_6;
  reg [31:0] coeffs_7;
  reg [31:0] coeffs_8;
  reg [31:0] coeffs_9;
  reg [31:0] coeffs_10;
  reg [31:0] coeffs_11;
  reg [31:0] coeffs_12;
  reg [31:0] coeffs_13;
  reg [31:0] coeffs_14;
  reg [31:0] coeffs_15;
  reg [31:0] coeffs_16;
  reg [31:0] coeffs_17;
  reg [31:0] coeffs_18;
  reg [31:0] coeffs_19;
  reg [31:0] coeffs_20;
  reg [31:0] coeffs_21;
  reg [31:0] coeffs_22;
  reg [31:0] coeffs_23;
  reg [31:0] coeffs_24;
  reg [31:0] coeffs_25;
  reg [31:0] coeffs_26;
  reg [31:0] coeffs_27;
  reg [31:0] coeffs_28;
  reg [31:0] coeffs_29;
  reg [31:0] coeffs_30;
  reg [31:0] coeffs_31;
  reg [31:0] coeffs_32;
  reg [31:0] coeffs_33;
  reg [31:0] coeffs_34;
  reg [31:0] coeffs_35;
  reg [31:0] coeffs_36;
  reg [31:0] coeffs_37;
  reg [31:0] coeffs_38;
  reg [31:0] coeffs_39;
  reg [31:0] coeffs_40;
  reg [31:0] coeffs_41;
  reg [31:0] coeffs_42;
  reg [31:0] coeffs_43;
  reg [31:0] coeffs_44;
  reg [31:0] coeffs_45;
  reg [31:0] coeffs_46;
  reg [31:0] coeffs_47;
  reg [31:0] coeffs_48;
  reg [31:0] coeffs_49;
  reg [31:0] coeffs_50;
  reg [31:0] coeffs_51;
  reg [31:0] coeffs_52;
  reg [31:0] coeffs_53;
  reg [31:0] coeffs_54;
  reg [31:0] coeffs_55;
  reg [31:0] coeffs_56;
  reg [31:0] coeffs_57;
  reg [31:0] coeffs_58;
  reg [31:0] coeffs_59;
  reg [31:0] coeffs_60;
  reg [31:0] coeffs_61;
  reg [31:0] coeffs_62;
  reg [31:0] coeffs_63;
  reg [31:0] coeffs_64;
  reg [31:0] coeffs_65;
  reg [31:0] coeffs_66;
  reg [31:0] coeffs_67;
  reg [31:0] coeffs_68;
  reg [31:0] coeffs_69;
  reg [31:0] coeffs_70;
  reg [31:0] coeffs_71;
  reg [31:0] coeffs_72;
  reg [31:0] coeffs_73;
  reg [31:0] coeffs_74;
  reg [31:0] coeffs_75;
  reg [31:0] coeffs_76;
  reg [31:0] coeffs_77;
  reg [31:0] coeffs_78;
  reg [31:0] coeffs_79;
  reg [31:0] coeffs_80;
  reg [31:0] coeffs_81;
  reg [31:0] coeffs_82;
  reg [31:0] coeffs_83;
  reg [31:0] coeffs_84;
  reg [31:0] coeffs_85;
  reg [31:0] coeffs_86;
  reg [31:0] coeffs_87;
  reg [31:0] coeffs_88;
  reg [31:0] coeffs_89;
  reg [31:0] coeffs_90;
  reg [31:0] coeffs_91;
  reg [31:0] coeffs_92;
  reg [31:0] coeffs_93;
  reg [31:0] coeffs_94;
  reg [31:0] coeffs_95;
  reg [31:0] coeffs_96;
  reg [31:0] coeffs_97;
  reg [31:0] coeffs_98;
  reg [31:0] coeffs_99;
  reg [31:0] data_0;
  reg [31:0] data_1;
  reg [31:0] data_2;
  reg [31:0] data_3;
  reg [31:0] data_4;
  reg [31:0] data_5;
  reg [31:0] data_6;
  reg [31:0] data_7;
  reg [31:0] data_8;
  reg [31:0] data_9;
  reg [31:0] data_10;
  reg [31:0] data_11;
  reg [31:0] data_12;
  reg [31:0] data_13;
  reg [31:0] data_14;
  reg [31:0] data_15;
  reg [31:0] data_16;
  reg [31:0] data_17;
  reg [31:0] data_18;
  reg [31:0] data_19;
  reg [31:0] data_20;
  reg [31:0] data_21;
  reg [31:0] data_22;
  reg [31:0] data_23;
  reg [31:0] data_24;
  reg [31:0] data_25;
  reg [31:0] data_26;
  reg [31:0] data_27;
  reg [31:0] data_28;
  reg [31:0] data_29;
  reg [31:0] data_30;
  reg [31:0] data_31;
  reg [31:0] data_32;
  reg [31:0] data_33;
  reg [31:0] data_34;
  reg [31:0] data_35;
  reg [31:0] data_36;
  reg [31:0] data_37;
  reg [31:0] data_38;
  reg [31:0] data_39;
  reg [31:0] data_40;
  reg [31:0] data_41;
  reg [31:0] data_42;
  reg [31:0] data_43;
  reg [31:0] data_44;
  reg [31:0] data_45;
  reg [31:0] data_46;
  reg [31:0] data_47;
  reg [31:0] data_48;
  reg [31:0] data_49;
  reg [31:0] data_50;
  reg [31:0] data_51;
  reg [31:0] data_52;
  reg [31:0] data_53;
  reg [31:0] data_54;
  reg [31:0] data_55;
  reg [31:0] data_56;
  reg [31:0] data_57;
  reg [31:0] data_58;
  reg [31:0] data_59;
  reg [31:0] data_60;
  reg [31:0] data_61;
  reg [31:0] data_62;
  reg [31:0] data_63;
  reg [31:0] data_64;
  reg [31:0] data_65;
  reg [31:0] data_66;
  reg [31:0] data_67;
  reg [31:0] data_68;
  reg [31:0] data_69;
  reg [31:0] data_70;
  reg [31:0] data_71;
  reg [31:0] data_72;
  reg [31:0] data_73;
  reg [31:0] data_74;
  reg [31:0] data_75;
  reg [31:0] data_76;
  reg [31:0] data_77;
  reg [31:0] data_78;
  reg [31:0] data_79;
  reg [31:0] data_80;
  reg [31:0] data_81;
  reg [31:0] data_82;
  reg [31:0] data_83;
  reg [31:0] data_84;
  reg [31:0] data_85;
  reg [31:0] data_86;
  reg [31:0] data_87;
  reg [31:0] data_88;
  reg [31:0] data_89;
  reg [31:0] data_90;
  reg [31:0] data_91;
  reg [31:0] data_92;
  reg [31:0] data_93;
  reg [31:0] data_94;
  reg [31:0] data_95;
  reg [31:0] data_96;
  reg [31:0] data_97;
  reg [31:0] data_98;
  reg [31:0] data_99;
  reg [63:0] result;
  wire [31:0] _GEN_101 = 7'h1 == rs2[6:0] ? $signed(coeffs_1) : $signed(coeffs_0);
  wire [31:0] _GEN_102 = 7'h2 == rs2[6:0] ? $signed(coeffs_2) : $signed(_GEN_101);
  wire [31:0] _GEN_103 = 7'h3 == rs2[6:0] ? $signed(coeffs_3) : $signed(_GEN_102);
  wire [31:0] _GEN_104 = 7'h4 == rs2[6:0] ? $signed(coeffs_4) : $signed(_GEN_103);
  wire [31:0] _GEN_105 = 7'h5 == rs2[6:0] ? $signed(coeffs_5) : $signed(_GEN_104);
  wire [31:0] _GEN_106 = 7'h6 == rs2[6:0] ? $signed(coeffs_6) : $signed(_GEN_105);
  wire [31:0] _GEN_107 = 7'h7 == rs2[6:0] ? $signed(coeffs_7) : $signed(_GEN_106);
  wire [31:0] _GEN_108 = 7'h8 == rs2[6:0] ? $signed(coeffs_8) : $signed(_GEN_107);
  wire [31:0] _GEN_109 = 7'h9 == rs2[6:0] ? $signed(coeffs_9) : $signed(_GEN_108);
  wire [31:0] _GEN_110 = 7'ha == rs2[6:0] ? $signed(coeffs_10) : $signed(_GEN_109);
  wire [31:0] _GEN_111 = 7'hb == rs2[6:0] ? $signed(coeffs_11) : $signed(_GEN_110);
  wire [31:0] _GEN_112 = 7'hc == rs2[6:0] ? $signed(coeffs_12) : $signed(_GEN_111);
  wire [31:0] _GEN_113 = 7'hd == rs2[6:0] ? $signed(coeffs_13) : $signed(_GEN_112);
  wire [31:0] _GEN_114 = 7'he == rs2[6:0] ? $signed(coeffs_14) : $signed(_GEN_113);
  wire [31:0] _GEN_115 = 7'hf == rs2[6:0] ? $signed(coeffs_15) : $signed(_GEN_114);
  wire [31:0] _GEN_116 = 7'h10 == rs2[6:0] ? $signed(coeffs_16) : $signed(_GEN_115);
  wire [31:0] _GEN_117 = 7'h11 == rs2[6:0] ? $signed(coeffs_17) : $signed(_GEN_116);
  wire [31:0] _GEN_118 = 7'h12 == rs2[6:0] ? $signed(coeffs_18) : $signed(_GEN_117);
  wire [31:0] _GEN_119 = 7'h13 == rs2[6:0] ? $signed(coeffs_19) : $signed(_GEN_118);
  wire [31:0] _GEN_120 = 7'h14 == rs2[6:0] ? $signed(coeffs_20) : $signed(_GEN_119);
  wire [31:0] _GEN_121 = 7'h15 == rs2[6:0] ? $signed(coeffs_21) : $signed(_GEN_120);
  wire [31:0] _GEN_122 = 7'h16 == rs2[6:0] ? $signed(coeffs_22) : $signed(_GEN_121);
  wire [31:0] _GEN_123 = 7'h17 == rs2[6:0] ? $signed(coeffs_23) : $signed(_GEN_122);
  wire [31:0] _GEN_124 = 7'h18 == rs2[6:0] ? $signed(coeffs_24) : $signed(_GEN_123);
  wire [31:0] _GEN_125 = 7'h19 == rs2[6:0] ? $signed(coeffs_25) : $signed(_GEN_124);
  wire [31:0] _GEN_126 = 7'h1a == rs2[6:0] ? $signed(coeffs_26) : $signed(_GEN_125);
  wire [31:0] _GEN_127 = 7'h1b == rs2[6:0] ? $signed(coeffs_27) : $signed(_GEN_126);
  wire [31:0] _GEN_128 = 7'h1c == rs2[6:0] ? $signed(coeffs_28) : $signed(_GEN_127);
  wire [31:0] _GEN_129 = 7'h1d == rs2[6:0] ? $signed(coeffs_29) : $signed(_GEN_128);
  wire [31:0] _GEN_130 = 7'h1e == rs2[6:0] ? $signed(coeffs_30) : $signed(_GEN_129);
  wire [31:0] _GEN_131 = 7'h1f == rs2[6:0] ? $signed(coeffs_31) : $signed(_GEN_130);
  wire [31:0] _GEN_132 = 7'h20 == rs2[6:0] ? $signed(coeffs_32) : $signed(_GEN_131);
  wire [31:0] _GEN_133 = 7'h21 == rs2[6:0] ? $signed(coeffs_33) : $signed(_GEN_132);
  wire [31:0] _GEN_134 = 7'h22 == rs2[6:0] ? $signed(coeffs_34) : $signed(_GEN_133);
  wire [31:0] _GEN_135 = 7'h23 == rs2[6:0] ? $signed(coeffs_35) : $signed(_GEN_134);
  wire [31:0] _GEN_136 = 7'h24 == rs2[6:0] ? $signed(coeffs_36) : $signed(_GEN_135);
  wire [31:0] _GEN_137 = 7'h25 == rs2[6:0] ? $signed(coeffs_37) : $signed(_GEN_136);
  wire [31:0] _GEN_138 = 7'h26 == rs2[6:0] ? $signed(coeffs_38) : $signed(_GEN_137);
  wire [31:0] _GEN_139 = 7'h27 == rs2[6:0] ? $signed(coeffs_39) : $signed(_GEN_138);
  wire [31:0] _GEN_140 = 7'h28 == rs2[6:0] ? $signed(coeffs_40) : $signed(_GEN_139);
  wire [31:0] _GEN_141 = 7'h29 == rs2[6:0] ? $signed(coeffs_41) : $signed(_GEN_140);
  wire [31:0] _GEN_142 = 7'h2a == rs2[6:0] ? $signed(coeffs_42) : $signed(_GEN_141);
  wire [31:0] _GEN_143 = 7'h2b == rs2[6:0] ? $signed(coeffs_43) : $signed(_GEN_142);
  wire [31:0] _GEN_144 = 7'h2c == rs2[6:0] ? $signed(coeffs_44) : $signed(_GEN_143);
  wire [31:0] _GEN_145 = 7'h2d == rs2[6:0] ? $signed(coeffs_45) : $signed(_GEN_144);
  wire [31:0] _GEN_146 = 7'h2e == rs2[6:0] ? $signed(coeffs_46) : $signed(_GEN_145);
  wire [31:0] _GEN_147 = 7'h2f == rs2[6:0] ? $signed(coeffs_47) : $signed(_GEN_146);
  wire [31:0] _GEN_148 = 7'h30 == rs2[6:0] ? $signed(coeffs_48) : $signed(_GEN_147);
  wire [31:0] _GEN_149 = 7'h31 == rs2[6:0] ? $signed(coeffs_49) : $signed(_GEN_148);
  wire [31:0] _GEN_150 = 7'h32 == rs2[6:0] ? $signed(coeffs_50) : $signed(_GEN_149);
  wire [31:0] _GEN_151 = 7'h33 == rs2[6:0] ? $signed(coeffs_51) : $signed(_GEN_150);
  wire [31:0] _GEN_152 = 7'h34 == rs2[6:0] ? $signed(coeffs_52) : $signed(_GEN_151);
  wire [31:0] _GEN_153 = 7'h35 == rs2[6:0] ? $signed(coeffs_53) : $signed(_GEN_152);
  wire [31:0] _GEN_154 = 7'h36 == rs2[6:0] ? $signed(coeffs_54) : $signed(_GEN_153);
  wire [31:0] _GEN_155 = 7'h37 == rs2[6:0] ? $signed(coeffs_55) : $signed(_GEN_154);
  wire [31:0] _GEN_156 = 7'h38 == rs2[6:0] ? $signed(coeffs_56) : $signed(_GEN_155);
  wire [31:0] _GEN_157 = 7'h39 == rs2[6:0] ? $signed(coeffs_57) : $signed(_GEN_156);
  wire [31:0] _GEN_158 = 7'h3a == rs2[6:0] ? $signed(coeffs_58) : $signed(_GEN_157);
  wire [31:0] _GEN_159 = 7'h3b == rs2[6:0] ? $signed(coeffs_59) : $signed(_GEN_158);
  wire [31:0] _GEN_160 = 7'h3c == rs2[6:0] ? $signed(coeffs_60) : $signed(_GEN_159);
  wire [31:0] _GEN_161 = 7'h3d == rs2[6:0] ? $signed(coeffs_61) : $signed(_GEN_160);
  wire [31:0] _GEN_162 = 7'h3e == rs2[6:0] ? $signed(coeffs_62) : $signed(_GEN_161);
  wire [31:0] _GEN_163 = 7'h3f == rs2[6:0] ? $signed(coeffs_63) : $signed(_GEN_162);
  wire [31:0] _GEN_164 = 7'h40 == rs2[6:0] ? $signed(coeffs_64) : $signed(_GEN_163);
  wire [31:0] _GEN_165 = 7'h41 == rs2[6:0] ? $signed(coeffs_65) : $signed(_GEN_164);
  wire [31:0] _GEN_166 = 7'h42 == rs2[6:0] ? $signed(coeffs_66) : $signed(_GEN_165);
  wire [31:0] _GEN_167 = 7'h43 == rs2[6:0] ? $signed(coeffs_67) : $signed(_GEN_166);
  wire [31:0] _GEN_168 = 7'h44 == rs2[6:0] ? $signed(coeffs_68) : $signed(_GEN_167);
  wire [31:0] _GEN_169 = 7'h45 == rs2[6:0] ? $signed(coeffs_69) : $signed(_GEN_168);
  wire [31:0] _GEN_170 = 7'h46 == rs2[6:0] ? $signed(coeffs_70) : $signed(_GEN_169);
  wire [31:0] _GEN_171 = 7'h47 == rs2[6:0] ? $signed(coeffs_71) : $signed(_GEN_170);
  wire [31:0] _GEN_172 = 7'h48 == rs2[6:0] ? $signed(coeffs_72) : $signed(_GEN_171);
  wire [31:0] _GEN_173 = 7'h49 == rs2[6:0] ? $signed(coeffs_73) : $signed(_GEN_172);
  wire [31:0] _GEN_174 = 7'h4a == rs2[6:0] ? $signed(coeffs_74) : $signed(_GEN_173);
  wire [31:0] _GEN_175 = 7'h4b == rs2[6:0] ? $signed(coeffs_75) : $signed(_GEN_174);
  wire [31:0] _GEN_176 = 7'h4c == rs2[6:0] ? $signed(coeffs_76) : $signed(_GEN_175);
  wire [31:0] _GEN_177 = 7'h4d == rs2[6:0] ? $signed(coeffs_77) : $signed(_GEN_176);
  wire [31:0] _GEN_178 = 7'h4e == rs2[6:0] ? $signed(coeffs_78) : $signed(_GEN_177);
  wire [31:0] _GEN_179 = 7'h4f == rs2[6:0] ? $signed(coeffs_79) : $signed(_GEN_178);
  wire [31:0] _GEN_180 = 7'h50 == rs2[6:0] ? $signed(coeffs_80) : $signed(_GEN_179);
  wire [31:0] _GEN_181 = 7'h51 == rs2[6:0] ? $signed(coeffs_81) : $signed(_GEN_180);
  wire [31:0] _GEN_182 = 7'h52 == rs2[6:0] ? $signed(coeffs_82) : $signed(_GEN_181);
  wire [31:0] _GEN_183 = 7'h53 == rs2[6:0] ? $signed(coeffs_83) : $signed(_GEN_182);
  wire [31:0] _GEN_184 = 7'h54 == rs2[6:0] ? $signed(coeffs_84) : $signed(_GEN_183);
  wire [31:0] _GEN_185 = 7'h55 == rs2[6:0] ? $signed(coeffs_85) : $signed(_GEN_184);
  wire [31:0] _GEN_186 = 7'h56 == rs2[6:0] ? $signed(coeffs_86) : $signed(_GEN_185);
  wire [31:0] _GEN_187 = 7'h57 == rs2[6:0] ? $signed(coeffs_87) : $signed(_GEN_186);
  wire [31:0] _GEN_188 = 7'h58 == rs2[6:0] ? $signed(coeffs_88) : $signed(_GEN_187);
  wire [31:0] _GEN_189 = 7'h59 == rs2[6:0] ? $signed(coeffs_89) : $signed(_GEN_188);
  wire [31:0] _GEN_190 = 7'h5a == rs2[6:0] ? $signed(coeffs_90) : $signed(_GEN_189);
  wire [31:0] _GEN_191 = 7'h5b == rs2[6:0] ? $signed(coeffs_91) : $signed(_GEN_190);
  wire [31:0] _GEN_192 = 7'h5c == rs2[6:0] ? $signed(coeffs_92) : $signed(_GEN_191);
  wire [31:0] _GEN_193 = 7'h5d == rs2[6:0] ? $signed(coeffs_93) : $signed(_GEN_192);
  wire [31:0] _GEN_194 = 7'h5e == rs2[6:0] ? $signed(coeffs_94) : $signed(_GEN_193);
  wire [31:0] _GEN_195 = 7'h5f == rs2[6:0] ? $signed(coeffs_95) : $signed(_GEN_194);
  wire [31:0] _GEN_196 = 7'h60 == rs2[6:0] ? $signed(coeffs_96) : $signed(_GEN_195);
  wire [31:0] _GEN_197 = 7'h61 == rs2[6:0] ? $signed(coeffs_97) : $signed(_GEN_196);
  wire [31:0] _GEN_198 = 7'h62 == rs2[6:0] ? $signed(coeffs_98) : $signed(_GEN_197);
  wire [31:0] _GEN_199 = 7'h63 == rs2[6:0] ? $signed(coeffs_99) : $signed(_GEN_198);
  wire [63:0] _result_T_2 = $signed(data_0) * $signed(coeffs_0);
  wire [63:0] _result_T_3 = $signed(data_1) * $signed(coeffs_1);
  wire [63:0] _result_T_4 = $signed(data_2) * $signed(coeffs_2);
  wire [63:0] _result_T_5 = $signed(data_3) * $signed(coeffs_3);
  wire [63:0] _result_T_6 = $signed(data_4) * $signed(coeffs_4);
  wire [63:0] _result_T_7 = $signed(data_5) * $signed(coeffs_5);
  wire [63:0] _result_T_8 = $signed(data_6) * $signed(coeffs_6);
  wire [63:0] _result_T_9 = $signed(data_7) * $signed(coeffs_7);
  wire [63:0] _result_T_10 = $signed(data_8) * $signed(coeffs_8);
  wire [63:0] _result_T_11 = $signed(data_9) * $signed(coeffs_9);
  wire [63:0] _result_T_12 = $signed(data_10) * $signed(coeffs_10);
  wire [63:0] _result_T_13 = $signed(data_11) * $signed(coeffs_11);
  wire [63:0] _result_T_14 = $signed(data_12) * $signed(coeffs_12);
  wire [63:0] _result_T_15 = $signed(data_13) * $signed(coeffs_13);
  wire [63:0] _result_T_16 = $signed(data_14) * $signed(coeffs_14);
  wire [63:0] _result_T_17 = $signed(data_15) * $signed(coeffs_15);
  wire [63:0] _result_T_18 = $signed(data_16) * $signed(coeffs_16);
  wire [63:0] _result_T_19 = $signed(data_17) * $signed(coeffs_17);
  wire [63:0] _result_T_20 = $signed(data_18) * $signed(coeffs_18);
  wire [63:0] _result_T_21 = $signed(data_19) * $signed(coeffs_19);
  wire [63:0] _result_T_22 = $signed(data_20) * $signed(coeffs_20);
  wire [63:0] _result_T_23 = $signed(data_21) * $signed(coeffs_21);
  wire [63:0] _result_T_24 = $signed(data_22) * $signed(coeffs_22);
  wire [63:0] _result_T_25 = $signed(data_23) * $signed(coeffs_23);
  wire [63:0] _result_T_26 = $signed(data_24) * $signed(coeffs_24);
  wire [63:0] _result_T_27 = $signed(data_25) * $signed(coeffs_25);
  wire [63:0] _result_T_28 = $signed(data_26) * $signed(coeffs_26);
  wire [63:0] _result_T_29 = $signed(data_27) * $signed(coeffs_27);
  wire [63:0] _result_T_30 = $signed(data_28) * $signed(coeffs_28);
  wire [63:0] _result_T_31 = $signed(data_29) * $signed(coeffs_29);
  wire [63:0] _result_T_32 = $signed(data_30) * $signed(coeffs_30);
  wire [63:0] _result_T_33 = $signed(data_31) * $signed(coeffs_31);
  wire [63:0] _result_T_34 = $signed(data_32) * $signed(coeffs_32);
  wire [63:0] _result_T_35 = $signed(data_33) * $signed(coeffs_33);
  wire [63:0] _result_T_36 = $signed(data_34) * $signed(coeffs_34);
  wire [63:0] _result_T_37 = $signed(data_35) * $signed(coeffs_35);
  wire [63:0] _result_T_38 = $signed(data_36) * $signed(coeffs_36);
  wire [63:0] _result_T_39 = $signed(data_37) * $signed(coeffs_37);
  wire [63:0] _result_T_40 = $signed(data_38) * $signed(coeffs_38);
  wire [63:0] _result_T_41 = $signed(data_39) * $signed(coeffs_39);
  wire [63:0] _result_T_42 = $signed(data_40) * $signed(coeffs_40);
  wire [63:0] _result_T_43 = $signed(data_41) * $signed(coeffs_41);
  wire [63:0] _result_T_44 = $signed(data_42) * $signed(coeffs_42);
  wire [63:0] _result_T_45 = $signed(data_43) * $signed(coeffs_43);
  wire [63:0] _result_T_46 = $signed(data_44) * $signed(coeffs_44);
  wire [63:0] _result_T_47 = $signed(data_45) * $signed(coeffs_45);
  wire [63:0] _result_T_48 = $signed(data_46) * $signed(coeffs_46);
  wire [63:0] _result_T_49 = $signed(data_47) * $signed(coeffs_47);
  wire [63:0] _result_T_50 = $signed(data_48) * $signed(coeffs_48);
  wire [63:0] _result_T_51 = $signed(data_49) * $signed(coeffs_49);
  wire [63:0] _result_T_52 = $signed(data_50) * $signed(coeffs_50);
  wire [63:0] _result_T_53 = $signed(data_51) * $signed(coeffs_51);
  wire [63:0] _result_T_54 = $signed(data_52) * $signed(coeffs_52);
  wire [63:0] _result_T_55 = $signed(data_53) * $signed(coeffs_53);
  wire [63:0] _result_T_56 = $signed(data_54) * $signed(coeffs_54);
  wire [63:0] _result_T_57 = $signed(data_55) * $signed(coeffs_55);
  wire [63:0] _result_T_58 = $signed(data_56) * $signed(coeffs_56);
  wire [63:0] _result_T_59 = $signed(data_57) * $signed(coeffs_57);
  wire [63:0] _result_T_60 = $signed(data_58) * $signed(coeffs_58);
  wire [63:0] _result_T_61 = $signed(data_59) * $signed(coeffs_59);
  wire [63:0] _result_T_62 = $signed(data_60) * $signed(coeffs_60);
  wire [63:0] _result_T_63 = $signed(data_61) * $signed(coeffs_61);
  wire [63:0] _result_T_64 = $signed(data_62) * $signed(coeffs_62);
  wire [63:0] _result_T_65 = $signed(data_63) * $signed(coeffs_63);
  wire [63:0] _result_T_66 = $signed(data_64) * $signed(coeffs_64);
  wire [63:0] _result_T_67 = $signed(data_65) * $signed(coeffs_65);
  wire [63:0] _result_T_68 = $signed(data_66) * $signed(coeffs_66);
  wire [63:0] _result_T_69 = $signed(data_67) * $signed(coeffs_67);
  wire [63:0] _result_T_70 = $signed(data_68) * $signed(coeffs_68);
  wire [63:0] _result_T_71 = $signed(data_69) * $signed(coeffs_69);
  wire [63:0] _result_T_72 = $signed(data_70) * $signed(coeffs_70);
  wire [63:0] _result_T_73 = $signed(data_71) * $signed(coeffs_71);
  wire [63:0] _result_T_74 = $signed(data_72) * $signed(coeffs_72);
  wire [63:0] _result_T_75 = $signed(data_73) * $signed(coeffs_73);
  wire [63:0] _result_T_76 = $signed(data_74) * $signed(coeffs_74);
  wire [63:0] _result_T_77 = $signed(data_75) * $signed(coeffs_75);
  wire [63:0] _result_T_78 = $signed(data_76) * $signed(coeffs_76);
  wire [63:0] _result_T_79 = $signed(data_77) * $signed(coeffs_77);
  wire [63:0] _result_T_80 = $signed(data_78) * $signed(coeffs_78);
  wire [63:0] _result_T_81 = $signed(data_79) * $signed(coeffs_79);
  wire [63:0] _result_T_82 = $signed(data_80) * $signed(coeffs_80);
  wire [63:0] _result_T_83 = $signed(data_81) * $signed(coeffs_81);
  wire [63:0] _result_T_84 = $signed(data_82) * $signed(coeffs_82);
  wire [63:0] _result_T_85 = $signed(data_83) * $signed(coeffs_83);
  wire [63:0] _result_T_86 = $signed(data_84) * $signed(coeffs_84);
  wire [63:0] _result_T_87 = $signed(data_85) * $signed(coeffs_85);
  wire [63:0] _result_T_88 = $signed(data_86) * $signed(coeffs_86);
  wire [63:0] _result_T_89 = $signed(data_87) * $signed(coeffs_87);
  wire [63:0] _result_T_90 = $signed(data_88) * $signed(coeffs_88);
  wire [63:0] _result_T_91 = $signed(data_89) * $signed(coeffs_89);
  wire [63:0] _result_T_92 = $signed(data_90) * $signed(coeffs_90);
  wire [63:0] _result_T_93 = $signed(data_91) * $signed(coeffs_91);
  wire [63:0] _result_T_94 = $signed(data_92) * $signed(coeffs_92);
  wire [63:0] _result_T_95 = $signed(data_93) * $signed(coeffs_93);
  wire [63:0] _result_T_96 = $signed(data_94) * $signed(coeffs_94);
  wire [63:0] _result_T_97 = $signed(data_95) * $signed(coeffs_95);
  wire [63:0] _result_T_98 = $signed(data_96) * $signed(coeffs_96);
  wire [63:0] _result_T_99 = $signed(data_97) * $signed(coeffs_97);
  wire [63:0] _result_T_100 = $signed(data_98) * $signed(coeffs_98);
  wire [63:0] _result_T_101 = $signed(data_99) * $signed(coeffs_99);
  wire [63:0] _result_T_104 = $signed(_result_T_2) + $signed(_result_T_3);
  wire [63:0] _result_T_107 = $signed(_result_T_104) + $signed(_result_T_4);
  wire [63:0] _result_T_110 = $signed(_result_T_107) + $signed(_result_T_5);
  wire [63:0] _result_T_113 = $signed(_result_T_110) + $signed(_result_T_6);
  wire [63:0] _result_T_116 = $signed(_result_T_113) + $signed(_result_T_7);
  wire [63:0] _result_T_119 = $signed(_result_T_116) + $signed(_result_T_8);
  wire [63:0] _result_T_122 = $signed(_result_T_119) + $signed(_result_T_9);
  wire [63:0] _result_T_125 = $signed(_result_T_122) + $signed(_result_T_10);
  wire [63:0] _result_T_128 = $signed(_result_T_125) + $signed(_result_T_11);
  wire [63:0] _result_T_131 = $signed(_result_T_128) + $signed(_result_T_12);
  wire [63:0] _result_T_134 = $signed(_result_T_131) + $signed(_result_T_13);
  wire [63:0] _result_T_137 = $signed(_result_T_134) + $signed(_result_T_14);
  wire [63:0] _result_T_140 = $signed(_result_T_137) + $signed(_result_T_15);
  wire [63:0] _result_T_143 = $signed(_result_T_140) + $signed(_result_T_16);
  wire [63:0] _result_T_146 = $signed(_result_T_143) + $signed(_result_T_17);
  wire [63:0] _result_T_149 = $signed(_result_T_146) + $signed(_result_T_18);
  wire [63:0] _result_T_152 = $signed(_result_T_149) + $signed(_result_T_19);
  wire [63:0] _result_T_155 = $signed(_result_T_152) + $signed(_result_T_20);
  wire [63:0] _result_T_158 = $signed(_result_T_155) + $signed(_result_T_21);
  wire [63:0] _result_T_161 = $signed(_result_T_158) + $signed(_result_T_22);
  wire [63:0] _result_T_164 = $signed(_result_T_161) + $signed(_result_T_23);
  wire [63:0] _result_T_167 = $signed(_result_T_164) + $signed(_result_T_24);
  wire [63:0] _result_T_170 = $signed(_result_T_167) + $signed(_result_T_25);
  wire [63:0] _result_T_173 = $signed(_result_T_170) + $signed(_result_T_26);
  wire [63:0] _result_T_176 = $signed(_result_T_173) + $signed(_result_T_27);
  wire [63:0] _result_T_179 = $signed(_result_T_176) + $signed(_result_T_28);
  wire [63:0] _result_T_182 = $signed(_result_T_179) + $signed(_result_T_29);
  wire [63:0] _result_T_185 = $signed(_result_T_182) + $signed(_result_T_30);
  wire [63:0] _result_T_188 = $signed(_result_T_185) + $signed(_result_T_31);
  wire [63:0] _result_T_191 = $signed(_result_T_188) + $signed(_result_T_32);
  wire [63:0] _result_T_194 = $signed(_result_T_191) + $signed(_result_T_33);
  wire [63:0] _result_T_197 = $signed(_result_T_194) + $signed(_result_T_34);
  wire [63:0] _result_T_200 = $signed(_result_T_197) + $signed(_result_T_35);
  wire [63:0] _result_T_203 = $signed(_result_T_200) + $signed(_result_T_36);
  wire [63:0] _result_T_206 = $signed(_result_T_203) + $signed(_result_T_37);
  wire [63:0] _result_T_209 = $signed(_result_T_206) + $signed(_result_T_38);
  wire [63:0] _result_T_212 = $signed(_result_T_209) + $signed(_result_T_39);
  wire [63:0] _result_T_215 = $signed(_result_T_212) + $signed(_result_T_40);
  wire [63:0] _result_T_218 = $signed(_result_T_215) + $signed(_result_T_41);
  wire [63:0] _result_T_221 = $signed(_result_T_218) + $signed(_result_T_42);
  wire [63:0] _result_T_224 = $signed(_result_T_221) + $signed(_result_T_43);
  wire [63:0] _result_T_227 = $signed(_result_T_224) + $signed(_result_T_44);
  wire [63:0] _result_T_230 = $signed(_result_T_227) + $signed(_result_T_45);
  wire [63:0] _result_T_233 = $signed(_result_T_230) + $signed(_result_T_46);
  wire [63:0] _result_T_236 = $signed(_result_T_233) + $signed(_result_T_47);
  wire [63:0] _result_T_239 = $signed(_result_T_236) + $signed(_result_T_48);
  wire [63:0] _result_T_242 = $signed(_result_T_239) + $signed(_result_T_49);
  wire [63:0] _result_T_245 = $signed(_result_T_242) + $signed(_result_T_50);
  wire [63:0] _result_T_248 = $signed(_result_T_245) + $signed(_result_T_51);
  wire [63:0] _result_T_251 = $signed(_result_T_248) + $signed(_result_T_52);
  wire [63:0] _result_T_254 = $signed(_result_T_251) + $signed(_result_T_53);
  wire [63:0] _result_T_257 = $signed(_result_T_254) + $signed(_result_T_54);
  wire [63:0] _result_T_260 = $signed(_result_T_257) + $signed(_result_T_55);
  wire [63:0] _result_T_263 = $signed(_result_T_260) + $signed(_result_T_56);
  wire [63:0] _result_T_266 = $signed(_result_T_263) + $signed(_result_T_57);
  wire [63:0] _result_T_269 = $signed(_result_T_266) + $signed(_result_T_58);
  wire [63:0] _result_T_272 = $signed(_result_T_269) + $signed(_result_T_59);
  wire [63:0] _result_T_275 = $signed(_result_T_272) + $signed(_result_T_60);
  wire [63:0] _result_T_278 = $signed(_result_T_275) + $signed(_result_T_61);
  wire [63:0] _result_T_281 = $signed(_result_T_278) + $signed(_result_T_62);
  wire [63:0] _result_T_284 = $signed(_result_T_281) + $signed(_result_T_63);
  wire [63:0] _result_T_287 = $signed(_result_T_284) + $signed(_result_T_64);
  wire [63:0] _result_T_290 = $signed(_result_T_287) + $signed(_result_T_65);
  wire [63:0] _result_T_293 = $signed(_result_T_290) + $signed(_result_T_66);
  wire [63:0] _result_T_296 = $signed(_result_T_293) + $signed(_result_T_67);
  wire [63:0] _result_T_299 = $signed(_result_T_296) + $signed(_result_T_68);
  wire [63:0] _result_T_302 = $signed(_result_T_299) + $signed(_result_T_69);
  wire [63:0] _result_T_305 = $signed(_result_T_302) + $signed(_result_T_70);
  wire [63:0] _result_T_308 = $signed(_result_T_305) + $signed(_result_T_71);
  wire [63:0] _result_T_311 = $signed(_result_T_308) + $signed(_result_T_72);
  wire [63:0] _result_T_314 = $signed(_result_T_311) + $signed(_result_T_73);
  wire [63:0] _result_T_317 = $signed(_result_T_314) + $signed(_result_T_74);
  wire [63:0] _result_T_320 = $signed(_result_T_317) + $signed(_result_T_75);
  wire [63:0] _result_T_323 = $signed(_result_T_320) + $signed(_result_T_76);
  wire [63:0] _result_T_326 = $signed(_result_T_323) + $signed(_result_T_77);
  wire [63:0] _result_T_329 = $signed(_result_T_326) + $signed(_result_T_78);
  wire [63:0] _result_T_332 = $signed(_result_T_329) + $signed(_result_T_79);
  wire [63:0] _result_T_335 = $signed(_result_T_332) + $signed(_result_T_80);
  wire [63:0] _result_T_338 = $signed(_result_T_335) + $signed(_result_T_81);
  wire [63:0] _result_T_341 = $signed(_result_T_338) + $signed(_result_T_82);
  wire [63:0] _result_T_344 = $signed(_result_T_341) + $signed(_result_T_83);
  wire [63:0] _result_T_347 = $signed(_result_T_344) + $signed(_result_T_84);
  wire [63:0] _result_T_350 = $signed(_result_T_347) + $signed(_result_T_85);
  wire [63:0] _result_T_353 = $signed(_result_T_350) + $signed(_result_T_86);
  wire [63:0] _result_T_356 = $signed(_result_T_353) + $signed(_result_T_87);
  wire [63:0] _result_T_359 = $signed(_result_T_356) + $signed(_result_T_88);
  wire [63:0] _result_T_362 = $signed(_result_T_359) + $signed(_result_T_89);
  wire [63:0] _result_T_365 = $signed(_result_T_362) + $signed(_result_T_90);
  wire [63:0] _result_T_368 = $signed(_result_T_365) + $signed(_result_T_91);
  wire [63:0] _result_T_371 = $signed(_result_T_368) + $signed(_result_T_92);
  wire [63:0] _result_T_374 = $signed(_result_T_371) + $signed(_result_T_93);
  wire [63:0] _result_T_377 = $signed(_result_T_374) + $signed(_result_T_94);
  wire [63:0] _result_T_380 = $signed(_result_T_377) + $signed(_result_T_95);
  wire [63:0] _result_T_383 = $signed(_result_T_380) + $signed(_result_T_96);
  wire [63:0] _result_T_386 = $signed(_result_T_383) + $signed(_result_T_97);
  wire [63:0] _result_T_389 = $signed(_result_T_386) + $signed(_result_T_98);
  wire [63:0] _result_T_392 = $signed(_result_T_389) + $signed(_result_T_99);
  wire [63:0] _result_T_395 = $signed(_result_T_392) + $signed(_result_T_100);
  wire [63:0] _result_T_398 = $signed(_result_T_395) + $signed(_result_T_101);
  wire [63:0] _GEN_200 = insn[6:0] == 7'h3b ? $signed(_result_T_398) : $signed(result);
  assign rd = result[31:0];
  always @(posedge clock) begin
    if (reset) begin
      coeffs_0 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h0 == rs2[6:0]) begin
          coeffs_0 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_1 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h1 == rs2[6:0]) begin
          coeffs_1 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_2 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h2 == rs2[6:0]) begin
          coeffs_2 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_3 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h3 == rs2[6:0]) begin
          coeffs_3 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_4 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h4 == rs2[6:0]) begin
          coeffs_4 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_5 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h5 == rs2[6:0]) begin
          coeffs_5 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_6 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h6 == rs2[6:0]) begin
          coeffs_6 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_7 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h7 == rs2[6:0]) begin
          coeffs_7 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_8 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h8 == rs2[6:0]) begin
          coeffs_8 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_9 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h9 == rs2[6:0]) begin
          coeffs_9 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_10 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'ha == rs2[6:0]) begin
          coeffs_10 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_11 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'hb == rs2[6:0]) begin
          coeffs_11 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_12 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'hc == rs2[6:0]) begin
          coeffs_12 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_13 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'hd == rs2[6:0]) begin
          coeffs_13 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_14 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'he == rs2[6:0]) begin
          coeffs_14 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_15 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'hf == rs2[6:0]) begin
          coeffs_15 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_16 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h10 == rs2[6:0]) begin
          coeffs_16 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_17 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h11 == rs2[6:0]) begin
          coeffs_17 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_18 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h12 == rs2[6:0]) begin
          coeffs_18 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_19 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h13 == rs2[6:0]) begin
          coeffs_19 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_20 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h14 == rs2[6:0]) begin
          coeffs_20 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_21 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h15 == rs2[6:0]) begin
          coeffs_21 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_22 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h16 == rs2[6:0]) begin
          coeffs_22 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_23 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h17 == rs2[6:0]) begin
          coeffs_23 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_24 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h18 == rs2[6:0]) begin
          coeffs_24 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_25 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h19 == rs2[6:0]) begin
          coeffs_25 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_26 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h1a == rs2[6:0]) begin
          coeffs_26 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_27 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h1b == rs2[6:0]) begin
          coeffs_27 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_28 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h1c == rs2[6:0]) begin
          coeffs_28 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_29 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h1d == rs2[6:0]) begin
          coeffs_29 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_30 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h1e == rs2[6:0]) begin
          coeffs_30 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_31 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h1f == rs2[6:0]) begin
          coeffs_31 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_32 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h20 == rs2[6:0]) begin
          coeffs_32 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_33 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h21 == rs2[6:0]) begin
          coeffs_33 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_34 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h22 == rs2[6:0]) begin
          coeffs_34 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_35 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h23 == rs2[6:0]) begin
          coeffs_35 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_36 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h24 == rs2[6:0]) begin
          coeffs_36 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_37 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h25 == rs2[6:0]) begin
          coeffs_37 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_38 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h26 == rs2[6:0]) begin
          coeffs_38 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_39 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h27 == rs2[6:0]) begin
          coeffs_39 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_40 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h28 == rs2[6:0]) begin
          coeffs_40 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_41 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h29 == rs2[6:0]) begin
          coeffs_41 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_42 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h2a == rs2[6:0]) begin
          coeffs_42 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_43 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h2b == rs2[6:0]) begin
          coeffs_43 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_44 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h2c == rs2[6:0]) begin
          coeffs_44 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_45 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h2d == rs2[6:0]) begin
          coeffs_45 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_46 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h2e == rs2[6:0]) begin
          coeffs_46 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_47 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h2f == rs2[6:0]) begin
          coeffs_47 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_48 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h30 == rs2[6:0]) begin
          coeffs_48 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_49 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h31 == rs2[6:0]) begin
          coeffs_49 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_50 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h32 == rs2[6:0]) begin
          coeffs_50 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_51 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h33 == rs2[6:0]) begin
          coeffs_51 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_52 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h34 == rs2[6:0]) begin
          coeffs_52 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_53 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h35 == rs2[6:0]) begin
          coeffs_53 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_54 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h36 == rs2[6:0]) begin
          coeffs_54 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_55 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h37 == rs2[6:0]) begin
          coeffs_55 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_56 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h38 == rs2[6:0]) begin
          coeffs_56 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_57 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h39 == rs2[6:0]) begin
          coeffs_57 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_58 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h3a == rs2[6:0]) begin
          coeffs_58 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_59 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h3b == rs2[6:0]) begin
          coeffs_59 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_60 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h3c == rs2[6:0]) begin
          coeffs_60 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_61 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h3d == rs2[6:0]) begin
          coeffs_61 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_62 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h3e == rs2[6:0]) begin
          coeffs_62 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_63 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h3f == rs2[6:0]) begin
          coeffs_63 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_64 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h40 == rs2[6:0]) begin
          coeffs_64 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_65 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h41 == rs2[6:0]) begin
          coeffs_65 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_66 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h42 == rs2[6:0]) begin
          coeffs_66 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_67 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h43 == rs2[6:0]) begin
          coeffs_67 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_68 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h44 == rs2[6:0]) begin
          coeffs_68 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_69 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h45 == rs2[6:0]) begin
          coeffs_69 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_70 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h46 == rs2[6:0]) begin
          coeffs_70 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_71 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h47 == rs2[6:0]) begin
          coeffs_71 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_72 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h48 == rs2[6:0]) begin
          coeffs_72 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_73 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h49 == rs2[6:0]) begin
          coeffs_73 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_74 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h4a == rs2[6:0]) begin
          coeffs_74 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_75 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h4b == rs2[6:0]) begin
          coeffs_75 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_76 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h4c == rs2[6:0]) begin
          coeffs_76 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_77 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h4d == rs2[6:0]) begin
          coeffs_77 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_78 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h4e == rs2[6:0]) begin
          coeffs_78 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_79 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h4f == rs2[6:0]) begin
          coeffs_79 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_80 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h50 == rs2[6:0]) begin
          coeffs_80 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_81 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h51 == rs2[6:0]) begin
          coeffs_81 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_82 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h52 == rs2[6:0]) begin
          coeffs_82 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_83 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h53 == rs2[6:0]) begin
          coeffs_83 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_84 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h54 == rs2[6:0]) begin
          coeffs_84 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_85 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h55 == rs2[6:0]) begin
          coeffs_85 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_86 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h56 == rs2[6:0]) begin
          coeffs_86 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_87 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h57 == rs2[6:0]) begin
          coeffs_87 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_88 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h58 == rs2[6:0]) begin
          coeffs_88 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_89 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h59 == rs2[6:0]) begin
          coeffs_89 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_90 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h5a == rs2[6:0]) begin
          coeffs_90 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_91 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h5b == rs2[6:0]) begin
          coeffs_91 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_92 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h5c == rs2[6:0]) begin
          coeffs_92 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_93 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h5d == rs2[6:0]) begin
          coeffs_93 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_94 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h5e == rs2[6:0]) begin
          coeffs_94 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_95 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h5f == rs2[6:0]) begin
          coeffs_95 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_96 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h60 == rs2[6:0]) begin
          coeffs_96 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_97 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h61 == rs2[6:0]) begin
          coeffs_97 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_98 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h62 == rs2[6:0]) begin
          coeffs_98 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_99 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h63 == rs2[6:0]) begin
          coeffs_99 <= rs1;
        end
      end
    end
    if (reset) begin
      data_0 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_0 <= rs1;
        end
      end
    end
    if (reset) begin
      data_1 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_1 <= data_0;
        end
      end
    end
    if (reset) begin
      data_2 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_2 <= data_1;
        end
      end
    end
    if (reset) begin
      data_3 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_3 <= data_2;
        end
      end
    end
    if (reset) begin
      data_4 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_4 <= data_3;
        end
      end
    end
    if (reset) begin
      data_5 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_5 <= data_4;
        end
      end
    end
    if (reset) begin
      data_6 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_6 <= data_5;
        end
      end
    end
    if (reset) begin
      data_7 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_7 <= data_6;
        end
      end
    end
    if (reset) begin
      data_8 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_8 <= data_7;
        end
      end
    end
    if (reset) begin
      data_9 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_9 <= data_8;
        end
      end
    end
    if (reset) begin
      data_10 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_10 <= data_9;
        end
      end
    end
    if (reset) begin
      data_11 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_11 <= data_10;
        end
      end
    end
    if (reset) begin
      data_12 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_12 <= data_11;
        end
      end
    end
    if (reset) begin
      data_13 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_13 <= data_12;
        end
      end
    end
    if (reset) begin
      data_14 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_14 <= data_13;
        end
      end
    end
    if (reset) begin
      data_15 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_15 <= data_14;
        end
      end
    end
    if (reset) begin
      data_16 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_16 <= data_15;
        end
      end
    end
    if (reset) begin
      data_17 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_17 <= data_16;
        end
      end
    end
    if (reset) begin
      data_18 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_18 <= data_17;
        end
      end
    end
    if (reset) begin
      data_19 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_19 <= data_18;
        end
      end
    end
    if (reset) begin
      data_20 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_20 <= data_19;
        end
      end
    end
    if (reset) begin
      data_21 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_21 <= data_20;
        end
      end
    end
    if (reset) begin
      data_22 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_22 <= data_21;
        end
      end
    end
    if (reset) begin
      data_23 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_23 <= data_22;
        end
      end
    end
    if (reset) begin
      data_24 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_24 <= data_23;
        end
      end
    end
    if (reset) begin
      data_25 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_25 <= data_24;
        end
      end
    end
    if (reset) begin
      data_26 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_26 <= data_25;
        end
      end
    end
    if (reset) begin
      data_27 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_27 <= data_26;
        end
      end
    end
    if (reset) begin
      data_28 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_28 <= data_27;
        end
      end
    end
    if (reset) begin
      data_29 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_29 <= data_28;
        end
      end
    end
    if (reset) begin
      data_30 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_30 <= data_29;
        end
      end
    end
    if (reset) begin
      data_31 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_31 <= data_30;
        end
      end
    end
    if (reset) begin
      data_32 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_32 <= data_31;
        end
      end
    end
    if (reset) begin
      data_33 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_33 <= data_32;
        end
      end
    end
    if (reset) begin
      data_34 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_34 <= data_33;
        end
      end
    end
    if (reset) begin
      data_35 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_35 <= data_34;
        end
      end
    end
    if (reset) begin
      data_36 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_36 <= data_35;
        end
      end
    end
    if (reset) begin
      data_37 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_37 <= data_36;
        end
      end
    end
    if (reset) begin
      data_38 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_38 <= data_37;
        end
      end
    end
    if (reset) begin
      data_39 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_39 <= data_38;
        end
      end
    end
    if (reset) begin
      data_40 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_40 <= data_39;
        end
      end
    end
    if (reset) begin
      data_41 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_41 <= data_40;
        end
      end
    end
    if (reset) begin
      data_42 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_42 <= data_41;
        end
      end
    end
    if (reset) begin
      data_43 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_43 <= data_42;
        end
      end
    end
    if (reset) begin
      data_44 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_44 <= data_43;
        end
      end
    end
    if (reset) begin
      data_45 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_45 <= data_44;
        end
      end
    end
    if (reset) begin
      data_46 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_46 <= data_45;
        end
      end
    end
    if (reset) begin
      data_47 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_47 <= data_46;
        end
      end
    end
    if (reset) begin
      data_48 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_48 <= data_47;
        end
      end
    end
    if (reset) begin
      data_49 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_49 <= data_48;
        end
      end
    end
    if (reset) begin
      data_50 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_50 <= data_49;
        end
      end
    end
    if (reset) begin
      data_51 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_51 <= data_50;
        end
      end
    end
    if (reset) begin
      data_52 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_52 <= data_51;
        end
      end
    end
    if (reset) begin
      data_53 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_53 <= data_52;
        end
      end
    end
    if (reset) begin
      data_54 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_54 <= data_53;
        end
      end
    end
    if (reset) begin
      data_55 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_55 <= data_54;
        end
      end
    end
    if (reset) begin
      data_56 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_56 <= data_55;
        end
      end
    end
    if (reset) begin
      data_57 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_57 <= data_56;
        end
      end
    end
    if (reset) begin
      data_58 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_58 <= data_57;
        end
      end
    end
    if (reset) begin
      data_59 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_59 <= data_58;
        end
      end
    end
    if (reset) begin
      data_60 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_60 <= data_59;
        end
      end
    end
    if (reset) begin
      data_61 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_61 <= data_60;
        end
      end
    end
    if (reset) begin
      data_62 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_62 <= data_61;
        end
      end
    end
    if (reset) begin
      data_63 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_63 <= data_62;
        end
      end
    end
    if (reset) begin
      data_64 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_64 <= data_63;
        end
      end
    end
    if (reset) begin
      data_65 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_65 <= data_64;
        end
      end
    end
    if (reset) begin
      data_66 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_66 <= data_65;
        end
      end
    end
    if (reset) begin
      data_67 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_67 <= data_66;
        end
      end
    end
    if (reset) begin
      data_68 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_68 <= data_67;
        end
      end
    end
    if (reset) begin
      data_69 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_69 <= data_68;
        end
      end
    end
    if (reset) begin
      data_70 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_70 <= data_69;
        end
      end
    end
    if (reset) begin
      data_71 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_71 <= data_70;
        end
      end
    end
    if (reset) begin
      data_72 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_72 <= data_71;
        end
      end
    end
    if (reset) begin
      data_73 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_73 <= data_72;
        end
      end
    end
    if (reset) begin
      data_74 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_74 <= data_73;
        end
      end
    end
    if (reset) begin
      data_75 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_75 <= data_74;
        end
      end
    end
    if (reset) begin
      data_76 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_76 <= data_75;
        end
      end
    end
    if (reset) begin
      data_77 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_77 <= data_76;
        end
      end
    end
    if (reset) begin
      data_78 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_78 <= data_77;
        end
      end
    end
    if (reset) begin
      data_79 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_79 <= data_78;
        end
      end
    end
    if (reset) begin
      data_80 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_80 <= data_79;
        end
      end
    end
    if (reset) begin
      data_81 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_81 <= data_80;
        end
      end
    end
    if (reset) begin
      data_82 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_82 <= data_81;
        end
      end
    end
    if (reset) begin
      data_83 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_83 <= data_82;
        end
      end
    end
    if (reset) begin
      data_84 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_84 <= data_83;
        end
      end
    end
    if (reset) begin
      data_85 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_85 <= data_84;
        end
      end
    end
    if (reset) begin
      data_86 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_86 <= data_85;
        end
      end
    end
    if (reset) begin
      data_87 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_87 <= data_86;
        end
      end
    end
    if (reset) begin
      data_88 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_88 <= data_87;
        end
      end
    end
    if (reset) begin
      data_89 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_89 <= data_88;
        end
      end
    end
    if (reset) begin
      data_90 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_90 <= data_89;
        end
      end
    end
    if (reset) begin
      data_91 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_91 <= data_90;
        end
      end
    end
    if (reset) begin
      data_92 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_92 <= data_91;
        end
      end
    end
    if (reset) begin
      data_93 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_93 <= data_92;
        end
      end
    end
    if (reset) begin
      data_94 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_94 <= data_93;
        end
      end
    end
    if (reset) begin
      data_95 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_95 <= data_94;
        end
      end
    end
    if (reset) begin
      data_96 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_96 <= data_95;
        end
      end
    end
    if (reset) begin
      data_97 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_97 <= data_96;
        end
      end
    end
    if (reset) begin
      data_98 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_98 <= data_97;
        end
      end
    end
    if (reset) begin
      data_99 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_99 <= data_98;
        end
      end
    end
    if (reset) begin
      result <= 64'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        result <= {{32{_GEN_199[31]}},_GEN_199};
      end else if (insn[6:0] == 7'h2b) begin
        result <= {{32{data_0[31]}},data_0};
      end else begin
        result <= _GEN_200;
      end
    end
  end
endmodule
