// SPDX-License-Identifier: Apache-2.0
// Example VCS Command: $VCS_HOME/bin/vcs -debug_pp -full64 +define+UNIT_DELAY +rad +v2k +vcs+lic+wait +vc+list +vcs+initreg+random +vcs+dumpvars+out.vcd tb.v SCIEPipelined.v ...
`timescale 100ps / 10ps

`define CLK_PERIOD 1

`define HALF_CLK_PERIOD 0.5
`define RESET_TIME 5
`define INIT_TIME 5.5
`define expect(nodeName, nodeVal, expVal, cycle) if (nodeVal !== expVal) begin \
  $display("\t ASSERTION ON %s FAILED @ CYCLE = %d, 0x%h != EXPECTED 0x%h", \
  nodeName,cycle,nodeVal,expVal); $stop; end

module testbench_v;

  integer cycle = 0;

  reg clock = 1;
  reg reset = 1;
  reg[31:0] io_rs2 = 0;
  reg signed [15:0] io_rs1_imag = 0;
  reg signed [15:0] io_rs1_real = 0;
  reg[31:0] io_insn = 0;
  reg[0:0] io_valid = 0;
  wire signed [15:0] io_rd_imag;
  wire signed [15:0] io_rd_real;

  always #`HALF_CLK_PERIOD clock = ~clock;

  initial begin
    #`RESET_TIME
    forever #`CLK_PERIOD cycle = cycle + 1;
  end

  SCIEPipelined SCIEPipelined(
    .clock(clock),
    .reset(reset),
    .io_rs2(io_rs2),
    .io_rs1_imag(io_rs1_imag),
    .io_rs1_real(io_rs1_real),
    .io_insn(io_insn),
    .io_valid(io_valid),
    .io_rd_imag(io_rd_imag),
    .io_rd_real(io_rd_real));

  initial begin
    #`INIT_TIME reset = 0;
    io_valid = 1'd1;
    io_insn = 4'd11;
    io_rs1_real = 5'd16;
    io_rs1_imag = -29;
    io_rs2 = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 4'd11;
    io_rs1_real = 5'd29;
    io_rs1_imag = -31;
    io_rs2 = 1'd1;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 4'd11;
    io_rs1_real = 6'd44;
    io_rs1_imag = -10;
    io_rs2 = 2'd2;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 4'd11;
    io_rs1_real = -17;
    io_rs1_imag = -18;
    io_rs2 = 2'd3;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 4'd11;
    io_rs1_real = -18;
    io_rs1_imag = -36;
    io_rs2 = 3'd4;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -47;
    io_rs1_imag = -48;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-2144,cycle)
    `expect("io_rd_imag",io_rd_imag,595,cycle)
    `expect("io_rd_real",io_rd_real,-2144,cycle)
    `expect("io_rd_imag",io_rd_imag,595,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -5;
    io_rs1_imag = 6'd40;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1771,cycle)
    `expect("io_rd_imag",io_rd_imag,850,cycle)
    `expect("io_rd_real",io_rd_real,-1771,cycle)
    `expect("io_rd_imag",io_rd_imag,850,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -29;
    io_rs1_imag = 5'd21;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1308,cycle)
    `expect("io_rd_imag",io_rd_imag,850,cycle)
    `expect("io_rd_real",io_rd_real,-1308,cycle)
    `expect("io_rd_imag",io_rd_imag,850,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -24;
    io_rs1_imag = 6'd32;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,469,cycle)
    `expect("io_rd_imag",io_rd_imag,6188,cycle)
    `expect("io_rd_real",io_rd_real,469,cycle)
    `expect("io_rd_imag",io_rd_imag,6188,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -44;
    io_rs1_imag = 3'd4;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1435,cycle)
    `expect("io_rd_imag",io_rd_imag,6192,cycle)
    `expect("io_rd_real",io_rd_real,-1435,cycle)
    `expect("io_rd_imag",io_rd_imag,6192,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 3'd5;
    io_rs1_imag = -11;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,274,cycle)
    `expect("io_rd_imag",io_rd_imag,2432,cycle)
    `expect("io_rd_real",io_rd_real,274,cycle)
    `expect("io_rd_imag",io_rd_imag,2432,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -29;
    io_rs1_imag = -28;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1106,cycle)
    `expect("io_rd_imag",io_rd_imag,1089,cycle)
    `expect("io_rd_real",io_rd_real,-1106,cycle)
    `expect("io_rd_imag",io_rd_imag,1089,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd38;
    io_rs1_imag = 2'd3;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1500,cycle)
    `expect("io_rd_imag",io_rd_imag,-489,cycle)
    `expect("io_rd_real",io_rd_real,1500,cycle)
    `expect("io_rd_imag",io_rd_imag,-489,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd40;
    io_rs1_imag = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,932,cycle)
    `expect("io_rd_imag",io_rd_imag,-1584,cycle)
    `expect("io_rd_real",io_rd_real,932,cycle)
    `expect("io_rd_imag",io_rd_imag,-1584,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -8;
    io_rs1_imag = -31;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1338,cycle)
    `expect("io_rd_imag",io_rd_imag,-736,cycle)
    `expect("io_rd_real",io_rd_real,1338,cycle)
    `expect("io_rd_imag",io_rd_imag,-736,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -19;
    io_rs1_imag = -17;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1308,cycle)
    `expect("io_rd_imag",io_rd_imag,41,cycle)
    `expect("io_rd_real",io_rd_real,-1308,cycle)
    `expect("io_rd_imag",io_rd_imag,41,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 3'd5;
    io_rs1_imag = -1;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-2945,cycle)
    `expect("io_rd_imag",io_rd_imag,-3491,cycle)
    `expect("io_rd_real",io_rd_real,-2945,cycle)
    `expect("io_rd_imag",io_rd_imag,-3491,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 4'd13;
    io_rs1_imag = -40;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-2986,cycle)
    `expect("io_rd_imag",io_rd_imag,-2528,cycle)
    `expect("io_rd_real",io_rd_real,-2986,cycle)
    `expect("io_rd_imag",io_rd_imag,-2528,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd36;
    io_rs1_imag = -23;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1699,cycle)
    `expect("io_rd_imag",io_rd_imag,-1592,cycle)
    `expect("io_rd_real",io_rd_real,-1699,cycle)
    `expect("io_rd_imag",io_rd_imag,-1592,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -11;
    io_rs1_imag = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-46,cycle)
    `expect("io_rd_imag",io_rd_imag,-2437,cycle)
    `expect("io_rd_real",io_rd_real,-46,cycle)
    `expect("io_rd_imag",io_rd_imag,-2437,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -8;
    io_rs1_imag = 5'd17;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,333,cycle)
    `expect("io_rd_imag",io_rd_imag,-243,cycle)
    `expect("io_rd_real",io_rd_real,333,cycle)
    `expect("io_rd_imag",io_rd_imag,-243,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd40;
    io_rs1_imag = 6'd37;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1176,cycle)
    `expect("io_rd_imag",io_rd_imag,278,cycle)
    `expect("io_rd_real",io_rd_real,-1176,cycle)
    `expect("io_rd_imag",io_rd_imag,278,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd27;
    io_rs1_imag = 6'd38;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,2370,cycle)
    `expect("io_rd_imag",io_rd_imag,-198,cycle)
    `expect("io_rd_real",io_rd_real,2370,cycle)
    `expect("io_rd_imag",io_rd_imag,-198,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd24;
    io_rs1_imag = -49;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,3694,cycle)
    `expect("io_rd_imag",io_rd_imag,264,cycle)
    `expect("io_rd_real",io_rd_real,3694,cycle)
    `expect("io_rd_imag",io_rd_imag,264,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -42;
    io_rs1_imag = -8;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,583,cycle)
    `expect("io_rd_imag",io_rd_imag,-1040,cycle)
    `expect("io_rd_real",io_rd_real,583,cycle)
    `expect("io_rd_imag",io_rd_imag,-1040,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd44;
    io_rs1_imag = 4'd10;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,931,cycle)
    `expect("io_rd_imag",io_rd_imag,-5680,cycle)
    `expect("io_rd_real",io_rd_real,931,cycle)
    `expect("io_rd_imag",io_rd_imag,-5680,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd24;
    io_rs1_imag = -1;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-395,cycle)
    `expect("io_rd_imag",io_rd_imag,-2973,cycle)
    `expect("io_rd_real",io_rd_real,-395,cycle)
    `expect("io_rd_imag",io_rd_imag,-2973,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 3'd5;
    io_rs1_imag = -21;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,546,cycle)
    `expect("io_rd_imag",io_rd_imag,-344,cycle)
    `expect("io_rd_real",io_rd_real,546,cycle)
    `expect("io_rd_imag",io_rd_imag,-344,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -40;
    io_rs1_imag = -41;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1389,cycle)
    `expect("io_rd_imag",io_rd_imag,150,cycle)
    `expect("io_rd_real",io_rd_real,-1389,cycle)
    `expect("io_rd_imag",io_rd_imag,150,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd46;
    io_rs1_imag = 6'd32;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1615,cycle)
    `expect("io_rd_imag",io_rd_imag,-3924,cycle)
    `expect("io_rd_real",io_rd_real,-1615,cycle)
    `expect("io_rd_imag",io_rd_imag,-3924,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -15;
    io_rs1_imag = -25;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1740,cycle)
    `expect("io_rd_imag",io_rd_imag,-2446,cycle)
    `expect("io_rd_real",io_rd_real,-1740,cycle)
    `expect("io_rd_imag",io_rd_imag,-2446,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -8;
    io_rs1_imag = 2'd2;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,160,cycle)
    `expect("io_rd_imag",io_rd_imag,2567,cycle)
    `expect("io_rd_real",io_rd_real,160,cycle)
    `expect("io_rd_imag",io_rd_imag,2567,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd46;
    io_rs1_imag = 2'd3;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1219,cycle)
    `expect("io_rd_imag",io_rd_imag,-1124,cycle)
    `expect("io_rd_real",io_rd_real,-1219,cycle)
    `expect("io_rd_imag",io_rd_imag,-1124,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd22;
    io_rs1_imag = -13;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1199,cycle)
    `expect("io_rd_imag",io_rd_imag,-3554,cycle)
    `expect("io_rd_real",io_rd_real,1199,cycle)
    `expect("io_rd_imag",io_rd_imag,-3554,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd43;
    io_rs1_imag = 3'd4;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,2635,cycle)
    `expect("io_rd_imag",io_rd_imag,-1470,cycle)
    `expect("io_rd_real",io_rd_real,2635,cycle)
    `expect("io_rd_imag",io_rd_imag,-1470,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 4'd10;
    io_rs1_imag = 6'd45;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,3162,cycle)
    `expect("io_rd_imag",io_rd_imag,-2206,cycle)
    `expect("io_rd_real",io_rd_real,3162,cycle)
    `expect("io_rd_imag",io_rd_imag,-2206,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -25;
    io_rs1_imag = -30;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1019,cycle)
    `expect("io_rd_imag",io_rd_imag,-899,cycle)
    `expect("io_rd_real",io_rd_real,1019,cycle)
    `expect("io_rd_imag",io_rd_imag,-899,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd33;
    io_rs1_imag = -22;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-2398,cycle)
    `expect("io_rd_imag",io_rd_imag,-924,cycle)
    `expect("io_rd_real",io_rd_real,-2398,cycle)
    `expect("io_rd_imag",io_rd_imag,-924,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -6;
    io_rs1_imag = -3;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1298,cycle)
    `expect("io_rd_imag",io_rd_imag,-5170,cycle)
    `expect("io_rd_real",io_rd_real,-1298,cycle)
    `expect("io_rd_imag",io_rd_imag,-5170,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -38;
    io_rs1_imag = -35;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,667,cycle)
    `expect("io_rd_imag",io_rd_imag,-867,cycle)
    `expect("io_rd_real",io_rd_real,667,cycle)
    `expect("io_rd_imag",io_rd_imag,-867,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -21;
    io_rs1_imag = 4'd8;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-4172,cycle)
    `expect("io_rd_imag",io_rd_imag,2048,cycle)
    `expect("io_rd_real",io_rd_real,-4172,cycle)
    `expect("io_rd_imag",io_rd_imag,2048,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd23;
    io_rs1_imag = 6'd34;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-2367,cycle)
    `expect("io_rd_imag",io_rd_imag,-1033,cycle)
    `expect("io_rd_real",io_rd_real,-2367,cycle)
    `expect("io_rd_imag",io_rd_imag,-1033,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd16;
    io_rs1_imag = -40;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-11,cycle)
    `expect("io_rd_imag",io_rd_imag,1280,cycle)
    `expect("io_rd_real",io_rd_real,-11,cycle)
    `expect("io_rd_imag",io_rd_imag,1280,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -13;
    io_rs1_imag = 5'd31;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1192,cycle)
    `expect("io_rd_imag",io_rd_imag,2723,cycle)
    `expect("io_rd_real",io_rd_real,1192,cycle)
    `expect("io_rd_imag",io_rd_imag,2723,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -38;
    io_rs1_imag = -42;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-51,cycle)
    `expect("io_rd_imag",io_rd_imag,-568,cycle)
    `expect("io_rd_real",io_rd_real,-51,cycle)
    `expect("io_rd_imag",io_rd_imag,-568,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 1'd0;
    io_rs1_imag = 2'd2;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-2790,cycle)
    `expect("io_rd_imag",io_rd_imag,438,cycle)
    `expect("io_rd_real",io_rd_real,-2790,cycle)
    `expect("io_rd_imag",io_rd_imag,438,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -35;
    io_rs1_imag = -12;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-3887,cycle)
    `expect("io_rd_imag",io_rd_imag,-736,cycle)
    `expect("io_rd_real",io_rd_real,-3887,cycle)
    `expect("io_rd_imag",io_rd_imag,-736,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -43;
    io_rs1_imag = -23;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1482,cycle)
    `expect("io_rd_imag",io_rd_imag,3012,cycle)
    `expect("io_rd_real",io_rd_real,-1482,cycle)
    `expect("io_rd_imag",io_rd_imag,3012,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd39;
    io_rs1_imag = -6;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-3962,cycle)
    `expect("io_rd_imag",io_rd_imag,1351,cycle)
    `expect("io_rd_real",io_rd_real,-3962,cycle)
    `expect("io_rd_imag",io_rd_imag,1351,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -16;
    io_rs1_imag = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-982,cycle)
    `expect("io_rd_imag",io_rd_imag,-703,cycle)
    `expect("io_rd_real",io_rd_real,-982,cycle)
    `expect("io_rd_imag",io_rd_imag,-703,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -47;
    io_rs1_imag = 6'd35;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1970,cycle)
    `expect("io_rd_imag",io_rd_imag,4406,cycle)
    `expect("io_rd_real",io_rd_real,1970,cycle)
    `expect("io_rd_imag",io_rd_imag,4406,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -37;
    io_rs1_imag = 3'd5;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-2254,cycle)
    `expect("io_rd_imag",io_rd_imag,5147,cycle)
    `expect("io_rd_real",io_rd_real,-2254,cycle)
    `expect("io_rd_imag",io_rd_imag,5147,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 1'd0;
    io_rs1_imag = -48;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-4674,cycle)
    `expect("io_rd_imag",io_rd_imag,1526,cycle)
    `expect("io_rd_real",io_rd_real,-4674,cycle)
    `expect("io_rd_imag",io_rd_imag,1526,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd32;
    io_rs1_imag = 4'd14;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-431,cycle)
    `expect("io_rd_imag",io_rd_imag,-679,cycle)
    `expect("io_rd_real",io_rd_real,-431,cycle)
    `expect("io_rd_imag",io_rd_imag,-679,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd46;
    io_rs1_imag = -24;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,3747,cycle)
    `expect("io_rd_imag",io_rd_imag,-2773,cycle)
    `expect("io_rd_real",io_rd_real,3747,cycle)
    `expect("io_rd_imag",io_rd_imag,-2773,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -5;
    io_rs1_imag = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,2040,cycle)
    `expect("io_rd_imag",io_rd_imag,377,cycle)
    `expect("io_rd_real",io_rd_real,2040,cycle)
    `expect("io_rd_imag",io_rd_imag,377,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -22;
    io_rs1_imag = 4'd11;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-414,cycle)
    `expect("io_rd_imag",io_rd_imag,-497,cycle)
    `expect("io_rd_real",io_rd_real,-414,cycle)
    `expect("io_rd_imag",io_rd_imag,-497,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -44;
    io_rs1_imag = -30;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-3377,cycle)
    `expect("io_rd_imag",io_rd_imag,23,cycle)
    `expect("io_rd_real",io_rd_real,-3377,cycle)
    `expect("io_rd_imag",io_rd_imag,23,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 3'd5;
    io_rs1_imag = -1;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-4620,cycle)
    `expect("io_rd_imag",io_rd_imag,-97,cycle)
    `expect("io_rd_real",io_rd_real,-4620,cycle)
    `expect("io_rd_imag",io_rd_imag,-97,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -9;
    io_rs1_imag = 5'd16;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1140,cycle)
    `expect("io_rd_imag",io_rd_imag,-158,cycle)
    `expect("io_rd_real",io_rd_real,-1140,cycle)
    `expect("io_rd_imag",io_rd_imag,-158,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -13;
    io_rs1_imag = -48;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-155,cycle)
    `expect("io_rd_imag",io_rd_imag,2154,cycle)
    `expect("io_rd_real",io_rd_real,-155,cycle)
    `expect("io_rd_imag",io_rd_imag,2154,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd45;
    io_rs1_imag = -30;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-2642,cycle)
    `expect("io_rd_imag",io_rd_imag,71,cycle)
    `expect("io_rd_real",io_rd_real,-2642,cycle)
    `expect("io_rd_imag",io_rd_imag,71,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -14;
    io_rs1_imag = -37;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1659,cycle)
    `expect("io_rd_imag",io_rd_imag,-4705,cycle)
    `expect("io_rd_real",io_rd_real,-1659,cycle)
    `expect("io_rd_imag",io_rd_imag,-4705,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -8;
    io_rs1_imag = -15;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-341,cycle)
    `expect("io_rd_imag",io_rd_imag,-1331,cycle)
    `expect("io_rd_real",io_rd_real,-341,cycle)
    `expect("io_rd_imag",io_rd_imag,-1331,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -6;
    io_rs1_imag = 6'd44;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-3302,cycle)
    `expect("io_rd_imag",io_rd_imag,235,cycle)
    `expect("io_rd_real",io_rd_real,-3302,cycle)
    `expect("io_rd_imag",io_rd_imag,235,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd26;
    io_rs1_imag = -16;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1678,cycle)
    `expect("io_rd_imag",io_rd_imag,-327,cycle)
    `expect("io_rd_real",io_rd_real,-1678,cycle)
    `expect("io_rd_imag",io_rd_imag,-327,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd18;
    io_rs1_imag = -22;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1130,cycle)
    `expect("io_rd_imag",io_rd_imag,1421,cycle)
    `expect("io_rd_real",io_rd_real,-1130,cycle)
    `expect("io_rd_imag",io_rd_imag,1421,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -21;
    io_rs1_imag = 5'd25;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1711,cycle)
    `expect("io_rd_imag",io_rd_imag,-1233,cycle)
    `expect("io_rd_real",io_rd_real,1711,cycle)
    `expect("io_rd_imag",io_rd_imag,-1233,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd46;
    io_rs1_imag = 6'd50;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,3886,cycle)
    `expect("io_rd_imag",io_rd_imag,-1078,cycle)
    `expect("io_rd_real",io_rd_real,3886,cycle)
    `expect("io_rd_imag",io_rd_imag,-1078,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 4'd13;
    io_rs1_imag = -37;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-401,cycle)
    `expect("io_rd_imag",io_rd_imag,-233,cycle)
    `expect("io_rd_real",io_rd_real,-401,cycle)
    `expect("io_rd_imag",io_rd_imag,-233,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd26;
    io_rs1_imag = -39;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,730,cycle)
    `expect("io_rd_imag",io_rd_imag,-1413,cycle)
    `expect("io_rd_real",io_rd_real,730,cycle)
    `expect("io_rd_imag",io_rd_imag,-1413,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 4'd9;
    io_rs1_imag = -1;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1258,cycle)
    `expect("io_rd_imag",io_rd_imag,-5344,cycle)
    `expect("io_rd_real",io_rd_real,1258,cycle)
    `expect("io_rd_imag",io_rd_imag,-5344,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -28;
    io_rs1_imag = 4'd11;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,940,cycle)
    `expect("io_rd_imag",io_rd_imag,-3457,cycle)
    `expect("io_rd_real",io_rd_real,940,cycle)
    `expect("io_rd_imag",io_rd_imag,-3457,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd29;
    io_rs1_imag = 6'd47;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-968,cycle)
    `expect("io_rd_imag",io_rd_imag,1357,cycle)
    `expect("io_rd_real",io_rd_real,-968,cycle)
    `expect("io_rd_imag",io_rd_imag,1357,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd27;
    io_rs1_imag = -25;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1160,cycle)
    `expect("io_rd_imag",io_rd_imag,-334,cycle)
    `expect("io_rd_real",io_rd_real,-1160,cycle)
    `expect("io_rd_imag",io_rd_imag,-334,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd44;
    io_rs1_imag = -25;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,2209,cycle)
    `expect("io_rd_imag",io_rd_imag,-1449,cycle)
    `expect("io_rd_real",io_rd_real,2209,cycle)
    `expect("io_rd_imag",io_rd_imag,-1449,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -8;
    io_rs1_imag = 4'd11;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,2883,cycle)
    `expect("io_rd_imag",io_rd_imag,-3562,cycle)
    `expect("io_rd_real",io_rd_real,2883,cycle)
    `expect("io_rd_imag",io_rd_imag,-3562,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 4'd10;
    io_rs1_imag = 6'd48;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,3608,cycle)
    `expect("io_rd_imag",io_rd_imag,-2446,cycle)
    `expect("io_rd_real",io_rd_real,3608,cycle)
    `expect("io_rd_imag",io_rd_imag,-2446,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd42;
    io_rs1_imag = -30;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1246,cycle)
    `expect("io_rd_imag",io_rd_imag,-941,cycle)
    `expect("io_rd_real",io_rd_real,-1246,cycle)
    `expect("io_rd_imag",io_rd_imag,-941,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -2;
    io_rs1_imag = 5'd20;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,398,cycle)
    `expect("io_rd_imag",io_rd_imag,-959,cycle)
    `expect("io_rd_real",io_rd_real,398,cycle)
    `expect("io_rd_imag",io_rd_imag,-959,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -23;
    io_rs1_imag = -33;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,2019,cycle)
    `expect("io_rd_imag",io_rd_imag,-1865,cycle)
    `expect("io_rd_real",io_rd_real,2019,cycle)
    `expect("io_rd_imag",io_rd_imag,-1865,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -22;
    io_rs1_imag = -5;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1781,cycle)
    `expect("io_rd_imag",io_rd_imag,-256,cycle)
    `expect("io_rd_real",io_rd_real,-1781,cycle)
    `expect("io_rd_imag",io_rd_imag,-256,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -38;
    io_rs1_imag = 6'd46;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-2851,cycle)
    `expect("io_rd_imag",io_rd_imag,-123,cycle)
    `expect("io_rd_real",io_rd_real,-2851,cycle)
    `expect("io_rd_imag",io_rd_imag,-123,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd42;
    io_rs1_imag = -20;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-49,cycle)
    `expect("io_rd_imag",io_rd_imag,1661,cycle)
    `expect("io_rd_real",io_rd_real,-49,cycle)
    `expect("io_rd_imag",io_rd_imag,1661,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd19;
    io_rs1_imag = 6'd41;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,389,cycle)
    `expect("io_rd_imag",io_rd_imag,2530,cycle)
    `expect("io_rd_real",io_rd_real,389,cycle)
    `expect("io_rd_imag",io_rd_imag,2530,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd48;
    io_rs1_imag = -13;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,5551,cycle)
    `expect("io_rd_imag",io_rd_imag,-1516,cycle)
    `expect("io_rd_real",io_rd_real,5551,cycle)
    `expect("io_rd_imag",io_rd_imag,-1516,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -14;
    io_rs1_imag = 5'd27;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,4060,cycle)
    `expect("io_rd_imag",io_rd_imag,711,cycle)
    `expect("io_rd_real",io_rd_real,4060,cycle)
    `expect("io_rd_imag",io_rd_imag,711,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd36;
    io_rs1_imag = 6'd43;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,3175,cycle)
    `expect("io_rd_imag",io_rd_imag,-2382,cycle)
    `expect("io_rd_real",io_rd_real,3175,cycle)
    `expect("io_rd_imag",io_rd_imag,-2382,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd25;
    io_rs1_imag = -40;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1355,cycle)
    `expect("io_rd_imag",io_rd_imag,-1971,cycle)
    `expect("io_rd_real",io_rd_real,1355,cycle)
    `expect("io_rd_imag",io_rd_imag,-1971,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd16;
    io_rs1_imag = -27;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,364,cycle)
    `expect("io_rd_imag",io_rd_imag,-3000,cycle)
    `expect("io_rd_real",io_rd_real,364,cycle)
    `expect("io_rd_imag",io_rd_imag,-3000,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -30;
    io_rs1_imag = -10;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,943,cycle)
    `expect("io_rd_imag",io_rd_imag,-3940,cycle)
    `expect("io_rd_real",io_rd_real,943,cycle)
    `expect("io_rd_imag",io_rd_imag,-3940,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -1;
    io_rs1_imag = -1;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1036,cycle)
    `expect("io_rd_imag",io_rd_imag,-2535,cycle)
    `expect("io_rd_real",io_rd_real,-1036,cycle)
    `expect("io_rd_imag",io_rd_imag,-2535,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd33;
    io_rs1_imag = 5'd30;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-2730,cycle)
    `expect("io_rd_imag",io_rd_imag,-624,cycle)
    `expect("io_rd_real",io_rd_real,-2730,cycle)
    `expect("io_rd_imag",io_rd_imag,-624,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 3'd4;
    io_rs1_imag = -13;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,590,cycle)
    `expect("io_rd_imag",io_rd_imag,109,cycle)
    `expect("io_rd_real",io_rd_real,590,cycle)
    `expect("io_rd_imag",io_rd_imag,109,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd31;
    io_rs1_imag = -4;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,2024,cycle)
    `expect("io_rd_imag",io_rd_imag,821,cycle)
    `expect("io_rd_real",io_rd_real,2024,cycle)
    `expect("io_rd_imag",io_rd_imag,821,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd42;
    io_rs1_imag = -23;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,787,cycle)
    `expect("io_rd_imag",io_rd_imag,-4325,cycle)
    `expect("io_rd_real",io_rd_real,787,cycle)
    `expect("io_rd_imag",io_rd_imag,-4325,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -16;
    io_rs1_imag = 5'd20;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,2337,cycle)
    `expect("io_rd_imag",io_rd_imag,-3250,cycle)
    `expect("io_rd_real",io_rd_real,2337,cycle)
    `expect("io_rd_imag",io_rd_imag,-3250,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -22;
    io_rs1_imag = 5'd20;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,863,cycle)
    `expect("io_rd_imag",io_rd_imag,202,cycle)
    `expect("io_rd_real",io_rd_real,863,cycle)
    `expect("io_rd_imag",io_rd_imag,202,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -26;
    io_rs1_imag = 6'd49;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1347,cycle)
    `expect("io_rd_imag",io_rd_imag,2431,cycle)
    `expect("io_rd_real",io_rd_real,-1347,cycle)
    `expect("io_rd_imag",io_rd_imag,2431,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -39;
    io_rs1_imag = -22;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-2217,cycle)
    `expect("io_rd_imag",io_rd_imag,2956,cycle)
    `expect("io_rd_real",io_rd_real,-2217,cycle)
    `expect("io_rd_imag",io_rd_imag,2956,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -15;
    io_rs1_imag = -8;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1197,cycle)
    `expect("io_rd_imag",io_rd_imag,3566,cycle)
    `expect("io_rd_real",io_rd_real,-1197,cycle)
    `expect("io_rd_imag",io_rd_imag,3566,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -35;
    io_rs1_imag = 4'd11;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-420,cycle)
    `expect("io_rd_imag",io_rd_imag,913,cycle)
    `expect("io_rd_real",io_rd_real,-420,cycle)
    `expect("io_rd_imag",io_rd_imag,913,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd23;
    io_rs1_imag = 5'd18;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1975,cycle)
    `expect("io_rd_imag",io_rd_imag,1953,cycle)
    `expect("io_rd_real",io_rd_real,1975,cycle)
    `expect("io_rd_imag",io_rd_imag,1953,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 4'd11;
    io_rs1_imag = 6'd43;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1239,cycle)
    `expect("io_rd_imag",io_rd_imag,3218,cycle)
    `expect("io_rd_real",io_rd_real,1239,cycle)
    `expect("io_rd_imag",io_rd_imag,3218,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd29;
    io_rs1_imag = 5'd19;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,4634,cycle)
    `expect("io_rd_imag",io_rd_imag,2058,cycle)
    `expect("io_rd_real",io_rd_real,4634,cycle)
    `expect("io_rd_imag",io_rd_imag,2058,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd42;
    io_rs1_imag = -5;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,3830,cycle)
    `expect("io_rd_imag",io_rd_imag,478,cycle)
    `expect("io_rd_real",io_rd_real,3830,cycle)
    `expect("io_rd_imag",io_rd_imag,478,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -37;
    io_rs1_imag = -41;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1569,cycle)
    `expect("io_rd_imag",io_rd_imag,-2565,cycle)
    `expect("io_rd_real",io_rd_real,1569,cycle)
    `expect("io_rd_imag",io_rd_imag,-2565,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 4'd15;
    io_rs1_imag = -31;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-6,cycle)
    `expect("io_rd_imag",io_rd_imag,-3628,cycle)
    `expect("io_rd_real",io_rd_real,-6,cycle)
    `expect("io_rd_imag",io_rd_imag,-3628,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 3'd5;
    io_rs1_imag = -5;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-3271,cycle)
    `expect("io_rd_imag",io_rd_imag,-5080,cycle)
    `expect("io_rd_real",io_rd_real,-3271,cycle)
    `expect("io_rd_imag",io_rd_imag,-5080,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 1'd1;
    io_rs1_imag = -19;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1240,cycle)
    `expect("io_rd_imag",io_rd_imag,-2206,cycle)
    `expect("io_rd_real",io_rd_real,-1240,cycle)
    `expect("io_rd_imag",io_rd_imag,-2206,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -9;
    io_rs1_imag = 5'd21;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1548,cycle)
    `expect("io_rd_imag",io_rd_imag,2072,cycle)
    `expect("io_rd_real",io_rd_real,-1548,cycle)
    `expect("io_rd_imag",io_rd_imag,2072,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd24;
    io_rs1_imag = 6'd48;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,459,cycle)
    `expect("io_rd_imag",io_rd_imag,127,cycle)
    `expect("io_rd_real",io_rd_real,459,cycle)
    `expect("io_rd_imag",io_rd_imag,127,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -15;
    io_rs1_imag = 6'd38;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,2231,cycle)
    `expect("io_rd_imag",io_rd_imag,2920,cycle)
    `expect("io_rd_real",io_rd_real,2231,cycle)
    `expect("io_rd_imag",io_rd_imag,2920,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -9;
    io_rs1_imag = -15;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1529,cycle)
    `expect("io_rd_imag",io_rd_imag,3571,cycle)
    `expect("io_rd_real",io_rd_real,1529,cycle)
    `expect("io_rd_imag",io_rd_imag,3571,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd32;
    io_rs1_imag = -28;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,68,cycle)
    `expect("io_rd_imag",io_rd_imag,-1012,cycle)
    `expect("io_rd_real",io_rd_real,68,cycle)
    `expect("io_rd_imag",io_rd_imag,-1012,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd31;
    io_rs1_imag = -33;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1288,cycle)
    `expect("io_rd_imag",io_rd_imag,-5905,cycle)
    `expect("io_rd_real",io_rd_real,1288,cycle)
    `expect("io_rd_imag",io_rd_imag,-5905,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd36;
    io_rs1_imag = -8;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,2869,cycle)
    `expect("io_rd_imag",io_rd_imag,-4369,cycle)
    `expect("io_rd_real",io_rd_real,2869,cycle)
    `expect("io_rd_imag",io_rd_imag,-4369,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd27;
    io_rs1_imag = 4'd14;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1242,cycle)
    `expect("io_rd_imag",io_rd_imag,-3175,cycle)
    `expect("io_rd_real",io_rd_real,1242,cycle)
    `expect("io_rd_imag",io_rd_imag,-3175,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd39;
    io_rs1_imag = 6'd42;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1858,cycle)
    `expect("io_rd_imag",io_rd_imag,-2247,cycle)
    `expect("io_rd_real",io_rd_real,1858,cycle)
    `expect("io_rd_imag",io_rd_imag,-2247,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 2'd2;
    io_rs1_imag = -2;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1233,cycle)
    `expect("io_rd_imag",io_rd_imag,-769,cycle)
    `expect("io_rd_real",io_rd_real,1233,cycle)
    `expect("io_rd_imag",io_rd_imag,-769,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -25;
    io_rs1_imag = 6'd40;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1749,cycle)
    `expect("io_rd_imag",io_rd_imag,827,cycle)
    `expect("io_rd_real",io_rd_real,1749,cycle)
    `expect("io_rd_imag",io_rd_imag,827,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd40;
    io_rs1_imag = 6'd34;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,2320,cycle)
    `expect("io_rd_imag",io_rd_imag,-1429,cycle)
    `expect("io_rd_real",io_rd_real,2320,cycle)
    `expect("io_rd_imag",io_rd_imag,-1429,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd48;
    io_rs1_imag = 2'd2;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,3080,cycle)
    `expect("io_rd_imag",io_rd_imag,-1766,cycle)
    `expect("io_rd_real",io_rd_real,3080,cycle)
    `expect("io_rd_imag",io_rd_imag,-1766,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -24;
    io_rs1_imag = -5;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,4062,cycle)
    `expect("io_rd_imag",io_rd_imag,16,cycle)
    `expect("io_rd_real",io_rd_real,4062,cycle)
    `expect("io_rd_imag",io_rd_imag,16,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -11;
    io_rs1_imag = 5'd27;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,3710,cycle)
    `expect("io_rd_imag",io_rd_imag,-160,cycle)
    `expect("io_rd_real",io_rd_real,3710,cycle)
    `expect("io_rd_imag",io_rd_imag,-160,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd26;
    io_rs1_imag = -44;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1724,cycle)
    `expect("io_rd_imag",io_rd_imag,-3264,cycle)
    `expect("io_rd_real",io_rd_real,-1724,cycle)
    `expect("io_rd_imag",io_rd_imag,-3264,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd37;
    io_rs1_imag = 3'd5;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-561,cycle)
    `expect("io_rd_imag",io_rd_imag,-3024,cycle)
    `expect("io_rd_real",io_rd_real,-561,cycle)
    `expect("io_rd_imag",io_rd_imag,-3024,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd41;
    io_rs1_imag = -38;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,2411,cycle)
    `expect("io_rd_imag",io_rd_imag,-4302,cycle)
    `expect("io_rd_real",io_rd_real,2411,cycle)
    `expect("io_rd_imag",io_rd_imag,-4302,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd46;
    io_rs1_imag = 5'd26;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,3115,cycle)
    `expect("io_rd_imag",io_rd_imag,-3251,cycle)
    `expect("io_rd_real",io_rd_real,3115,cycle)
    `expect("io_rd_imag",io_rd_imag,-3251,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -46;
    io_rs1_imag = 5'd16;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,701,cycle)
    `expect("io_rd_imag",io_rd_imag,-2059,cycle)
    `expect("io_rd_real",io_rd_real,701,cycle)
    `expect("io_rd_imag",io_rd_imag,-2059,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -42;
    io_rs1_imag = 5'd27;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-310,cycle)
    `expect("io_rd_imag",io_rd_imag,2710,cycle)
    `expect("io_rd_real",io_rd_real,-310,cycle)
    `expect("io_rd_imag",io_rd_imag,2710,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -39;
    io_rs1_imag = -48;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-6681,cycle)
    `expect("io_rd_imag",io_rd_imag,1550,cycle)
    `expect("io_rd_real",io_rd_real,-6681,cycle)
    `expect("io_rd_imag",io_rd_imag,1550,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -34;
    io_rs1_imag = -24;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-4259,cycle)
    `expect("io_rd_imag",io_rd_imag,459,cycle)
    `expect("io_rd_real",io_rd_real,-4259,cycle)
    `expect("io_rd_imag",io_rd_imag,459,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -40;
    io_rs1_imag = 5'd30;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1092,cycle)
    `expect("io_rd_imag",io_rd_imag,1941,cycle)
    `expect("io_rd_real",io_rd_real,-1092,cycle)
    `expect("io_rd_imag",io_rd_imag,1941,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 4'd8;
    io_rs1_imag = -1;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-340,cycle)
    `expect("io_rd_imag",io_rd_imag,3690,cycle)
    `expect("io_rd_real",io_rd_real,-340,cycle)
    `expect("io_rd_imag",io_rd_imag,3690,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -47;
    io_rs1_imag = -25;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-3616,cycle)
    `expect("io_rd_imag",io_rd_imag,5694,cycle)
    `expect("io_rd_real",io_rd_real,-3616,cycle)
    `expect("io_rd_imag",io_rd_imag,5694,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 1'd0;
    io_rs1_imag = 3'd6;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-654,cycle)
    `expect("io_rd_imag",io_rd_imag,2570,cycle)
    `expect("io_rd_real",io_rd_real,-654,cycle)
    `expect("io_rd_imag",io_rd_imag,2570,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -24;
    io_rs1_imag = -34;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1856,cycle)
    `expect("io_rd_imag",io_rd_imag,469,cycle)
    `expect("io_rd_real",io_rd_real,-1856,cycle)
    `expect("io_rd_imag",io_rd_imag,469,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -41;
    io_rs1_imag = 6'd42;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-959,cycle)
    `expect("io_rd_imag",io_rd_imag,2884,cycle)
    `expect("io_rd_real",io_rd_real,-959,cycle)
    `expect("io_rd_imag",io_rd_imag,2884,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -21;
    io_rs1_imag = -49;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-2986,cycle)
    `expect("io_rd_imag",io_rd_imag,3098,cycle)
    `expect("io_rd_real",io_rd_real,-2986,cycle)
    `expect("io_rd_imag",io_rd_imag,3098,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd45;
    io_rs1_imag = 6'd45;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1475,cycle)
    `expect("io_rd_imag",io_rd_imag,1805,cycle)
    `expect("io_rd_real",io_rd_real,-1475,cycle)
    `expect("io_rd_imag",io_rd_imag,1805,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -21;
    io_rs1_imag = 5'd21;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,2220,cycle)
    `expect("io_rd_imag",io_rd_imag,409,cycle)
    `expect("io_rd_real",io_rd_real,2220,cycle)
    `expect("io_rd_imag",io_rd_imag,409,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 4'd9;
    io_rs1_imag = -40;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,3181,cycle)
    `expect("io_rd_imag",io_rd_imag,3820,cycle)
    `expect("io_rd_real",io_rd_real,3181,cycle)
    `expect("io_rd_imag",io_rd_imag,3820,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -47;
    io_rs1_imag = -6;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-3960,cycle)
    `expect("io_rd_imag",io_rd_imag,1025,cycle)
    `expect("io_rd_real",io_rd_real,-3960,cycle)
    `expect("io_rd_imag",io_rd_imag,1025,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 2'd3;
    io_rs1_imag = 6'd43;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1287,cycle)
    `expect("io_rd_imag",io_rd_imag,-2375,cycle)
    `expect("io_rd_real",io_rd_real,1287,cycle)
    `expect("io_rd_imag",io_rd_imag,-2375,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -7;
    io_rs1_imag = -26;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1313,cycle)
    `expect("io_rd_imag",io_rd_imag,2043,cycle)
    `expect("io_rd_real",io_rd_real,-1313,cycle)
    `expect("io_rd_imag",io_rd_imag,2043,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd31;
    io_rs1_imag = -37;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1935,cycle)
    `expect("io_rd_imag",io_rd_imag,1178,cycle)
    `expect("io_rd_real",io_rd_real,-1935,cycle)
    `expect("io_rd_imag",io_rd_imag,1178,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 2'd2;
    io_rs1_imag = -36;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-475,cycle)
    `expect("io_rd_imag",io_rd_imag,-2727,cycle)
    `expect("io_rd_real",io_rd_real,-475,cycle)
    `expect("io_rd_imag",io_rd_imag,-2727,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 3'd5;
    io_rs1_imag = 4'd9;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1422,cycle)
    `expect("io_rd_imag",io_rd_imag,-3359,cycle)
    `expect("io_rd_real",io_rd_real,1422,cycle)
    `expect("io_rd_imag",io_rd_imag,-3359,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -6;
    io_rs1_imag = 3'd5;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1802,cycle)
    `expect("io_rd_imag",io_rd_imag,-453,cycle)
    `expect("io_rd_real",io_rd_real,-1802,cycle)
    `expect("io_rd_imag",io_rd_imag,-453,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 3'd5;
    io_rs1_imag = -3;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-2288,cycle)
    `expect("io_rd_imag",io_rd_imag,610,cycle)
    `expect("io_rd_real",io_rd_real,-2288,cycle)
    `expect("io_rd_imag",io_rd_imag,610,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -46;
    io_rs1_imag = -13;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-2530,cycle)
    `expect("io_rd_imag",io_rd_imag,1497,cycle)
    `expect("io_rd_real",io_rd_real,-2530,cycle)
    `expect("io_rd_imag",io_rd_imag,1497,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd39;
    io_rs1_imag = -14;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-903,cycle)
    `expect("io_rd_imag",io_rd_imag,-807,cycle)
    `expect("io_rd_real",io_rd_real,-903,cycle)
    `expect("io_rd_imag",io_rd_imag,-807,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -13;
    io_rs1_imag = -41;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-2705,cycle)
    `expect("io_rd_imag",io_rd_imag,-1919,cycle)
    `expect("io_rd_real",io_rd_real,-2705,cycle)
    `expect("io_rd_imag",io_rd_imag,-1919,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -41;
    io_rs1_imag = -19;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-929,cycle)
    `expect("io_rd_imag",io_rd_imag,16,cycle)
    `expect("io_rd_real",io_rd_real,-929,cycle)
    `expect("io_rd_imag",io_rd_imag,16,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd20;
    io_rs1_imag = -28;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-3807,cycle)
    `expect("io_rd_imag",io_rd_imag,-556,cycle)
    `expect("io_rd_real",io_rd_real,-3807,cycle)
    `expect("io_rd_imag",io_rd_imag,-556,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -20;
    io_rs1_imag = -19;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-4876,cycle)
    `expect("io_rd_imag",io_rd_imag,-1803,cycle)
    `expect("io_rd_real",io_rd_real,-4876,cycle)
    `expect("io_rd_imag",io_rd_imag,-1803,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -44;
    io_rs1_imag = -33;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-3117,cycle)
    `expect("io_rd_imag",io_rd_imag,1652,cycle)
    `expect("io_rd_real",io_rd_real,-3117,cycle)
    `expect("io_rd_imag",io_rd_imag,1652,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd44;
    io_rs1_imag = -30;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-4325,cycle)
    `expect("io_rd_imag",io_rd_imag,-51,cycle)
    `expect("io_rd_real",io_rd_real,-4325,cycle)
    `expect("io_rd_imag",io_rd_imag,-51,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd27;
    io_rs1_imag = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-2858,cycle)
    `expect("io_rd_imag",io_rd_imag,-3562,cycle)
    `expect("io_rd_real",io_rd_real,-2858,cycle)
    `expect("io_rd_imag",io_rd_imag,-3562,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -30;
    io_rs1_imag = 6'd47;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,3132,cycle)
    `expect("io_rd_imag",io_rd_imag,1440,cycle)
    `expect("io_rd_real",io_rd_real,3132,cycle)
    `expect("io_rd_imag",io_rd_imag,1440,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd33;
    io_rs1_imag = -29;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-222,cycle)
    `expect("io_rd_imag",io_rd_imag,2498,cycle)
    `expect("io_rd_real",io_rd_real,-222,cycle)
    `expect("io_rd_imag",io_rd_imag,2498,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 4'd11;
    io_rs1_imag = 6'd38;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1845,cycle)
    `expect("io_rd_imag",io_rd_imag,-737,cycle)
    `expect("io_rd_real",io_rd_real,-1845,cycle)
    `expect("io_rd_imag",io_rd_imag,-737,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 2'd3;
    io_rs1_imag = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,3577,cycle)
    `expect("io_rd_imag",io_rd_imag,-2163,cycle)
    `expect("io_rd_real",io_rd_real,3577,cycle)
    `expect("io_rd_imag",io_rd_imag,-2163,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd45;
    io_rs1_imag = 5'd18;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,3342,cycle)
    `expect("io_rd_imag",io_rd_imag,585,cycle)
    `expect("io_rd_real",io_rd_real,3342,cycle)
    `expect("io_rd_imag",io_rd_imag,585,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd18;
    io_rs1_imag = 5'd28;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1954,cycle)
    `expect("io_rd_imag",io_rd_imag,-2487,cycle)
    `expect("io_rd_real",io_rd_real,1954,cycle)
    `expect("io_rd_imag",io_rd_imag,-2487,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd26;
    io_rs1_imag = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,5085,cycle)
    `expect("io_rd_imag",io_rd_imag,-1292,cycle)
    `expect("io_rd_real",io_rd_real,5085,cycle)
    `expect("io_rd_imag",io_rd_imag,-1292,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -14;
    io_rs1_imag = -32;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,179,cycle)
    `expect("io_rd_imag",io_rd_imag,-1084,cycle)
    `expect("io_rd_real",io_rd_real,179,cycle)
    `expect("io_rd_imag",io_rd_imag,-1084,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd29;
    io_rs1_imag = 6'd43;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1493,cycle)
    `expect("io_rd_imag",io_rd_imag,-3651,cycle)
    `expect("io_rd_real",io_rd_real,1493,cycle)
    `expect("io_rd_imag",io_rd_imag,-3651,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd37;
    io_rs1_imag = -11;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1753,cycle)
    `expect("io_rd_imag",io_rd_imag,-3789,cycle)
    `expect("io_rd_real",io_rd_real,1753,cycle)
    `expect("io_rd_imag",io_rd_imag,-3789,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -44;
    io_rs1_imag = 5'd18;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1450,cycle)
    `expect("io_rd_imag",io_rd_imag,1560,cycle)
    `expect("io_rd_real",io_rd_real,1450,cycle)
    `expect("io_rd_imag",io_rd_imag,1560,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -15;
    io_rs1_imag = 2'd3;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,28,cycle)
    `expect("io_rd_imag",io_rd_imag,1342,cycle)
    `expect("io_rd_real",io_rd_real,28,cycle)
    `expect("io_rd_imag",io_rd_imag,1342,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd47;
    io_rs1_imag = -16;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1611,cycle)
    `expect("io_rd_imag",io_rd_imag,-2132,cycle)
    `expect("io_rd_real",io_rd_real,-1611,cycle)
    `expect("io_rd_imag",io_rd_imag,-2132,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -39;
    io_rs1_imag = -36;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1421,cycle)
    `expect("io_rd_imag",io_rd_imag,-1732,cycle)
    `expect("io_rd_real",io_rd_real,-1421,cycle)
    `expect("io_rd_imag",io_rd_imag,-1732,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -44;
    io_rs1_imag = 4'd15;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1141,cycle)
    `expect("io_rd_imag",io_rd_imag,1986,cycle)
    `expect("io_rd_real",io_rd_real,1141,cycle)
    `expect("io_rd_imag",io_rd_imag,1986,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -21;
    io_rs1_imag = 6'd40;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-2772,cycle)
    `expect("io_rd_imag",io_rd_imag,1766,cycle)
    `expect("io_rd_real",io_rd_real,-2772,cycle)
    `expect("io_rd_imag",io_rd_imag,1766,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd25;
    io_rs1_imag = -34;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-3148,cycle)
    `expect("io_rd_imag",io_rd_imag,1552,cycle)
    `expect("io_rd_real",io_rd_real,-3148,cycle)
    `expect("io_rd_imag",io_rd_imag,1552,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd17;
    io_rs1_imag = -38;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1259,cycle)
    `expect("io_rd_imag",io_rd_imag,1697,cycle)
    `expect("io_rd_real",io_rd_real,-1259,cycle)
    `expect("io_rd_imag",io_rd_imag,1697,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -2;
    io_rs1_imag = 5'd29;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,3293,cycle)
    `expect("io_rd_imag",io_rd_imag,-1841,cycle)
    `expect("io_rd_real",io_rd_real,3293,cycle)
    `expect("io_rd_imag",io_rd_imag,-1841,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd38;
    io_rs1_imag = -34;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1612,cycle)
    `expect("io_rd_imag",io_rd_imag,-2421,cycle)
    `expect("io_rd_real",io_rd_real,1612,cycle)
    `expect("io_rd_imag",io_rd_imag,-2421,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -45;
    io_rs1_imag = 6'd48;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1725,cycle)
    `expect("io_rd_imag",io_rd_imag,1257,cycle)
    `expect("io_rd_real",io_rd_real,-1725,cycle)
    `expect("io_rd_imag",io_rd_imag,1257,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd17;
    io_rs1_imag = -33;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-288,cycle)
    `expect("io_rd_imag",io_rd_imag,-495,cycle)
    `expect("io_rd_real",io_rd_real,-288,cycle)
    `expect("io_rd_imag",io_rd_imag,-495,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -45;
    io_rs1_imag = 3'd4;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-2812,cycle)
    `expect("io_rd_imag",io_rd_imag,1891,cycle)
    `expect("io_rd_real",io_rd_real,-2812,cycle)
    `expect("io_rd_imag",io_rd_imag,1891,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -9;
    io_rs1_imag = 6'd33;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-229,cycle)
    `expect("io_rd_imag",io_rd_imag,-84,cycle)
    `expect("io_rd_real",io_rd_real,-229,cycle)
    `expect("io_rd_imag",io_rd_imag,-84,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -38;
    io_rs1_imag = 5'd21;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,478,cycle)
    `expect("io_rd_imag",io_rd_imag,4311,cycle)
    `expect("io_rd_real",io_rd_real,478,cycle)
    `expect("io_rd_imag",io_rd_imag,4311,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd26;
    io_rs1_imag = -41;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1947,cycle)
    `expect("io_rd_imag",io_rd_imag,2643,cycle)
    `expect("io_rd_real",io_rd_real,-1947,cycle)
    `expect("io_rd_imag",io_rd_imag,2643,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd22;
    io_rs1_imag = 3'd5;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,219,cycle)
    `expect("io_rd_imag",io_rd_imag,-100,cycle)
    `expect("io_rd_real",io_rd_real,219,cycle)
    `expect("io_rd_imag",io_rd_imag,-100,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -4;
    io_rs1_imag = 4'd15;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,4272,cycle)
    `expect("io_rd_imag",io_rd_imag,-2188,cycle)
    `expect("io_rd_real",io_rd_real,4272,cycle)
    `expect("io_rd_imag",io_rd_imag,-2188,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd21;
    io_rs1_imag = 5'd22;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,2601,cycle)
    `expect("io_rd_imag",io_rd_imag,1521,cycle)
    `expect("io_rd_real",io_rd_real,2601,cycle)
    `expect("io_rd_imag",io_rd_imag,1521,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -23;
    io_rs1_imag = 6'd46;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,3,cycle)
    `expect("io_rd_imag",io_rd_imag,1411,cycle)
    `expect("io_rd_real",io_rd_real,3,cycle)
    `expect("io_rd_imag",io_rd_imag,1411,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd19;
    io_rs1_imag = 5'd23;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,2996,cycle)
    `expect("io_rd_imag",io_rd_imag,1557,cycle)
    `expect("io_rd_real",io_rd_real,2996,cycle)
    `expect("io_rd_imag",io_rd_imag,1557,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -15;
    io_rs1_imag = 5'd23;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1790,cycle)
    `expect("io_rd_imag",io_rd_imag,2257,cycle)
    `expect("io_rd_real",io_rd_real,1790,cycle)
    `expect("io_rd_imag",io_rd_imag,2257,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd44;
    io_rs1_imag = 1'd1;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,3710,cycle)
    `expect("io_rd_imag",io_rd_imag,-826,cycle)
    `expect("io_rd_real",io_rd_real,3710,cycle)
    `expect("io_rd_imag",io_rd_imag,-826,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 4'd11;
    io_rs1_imag = 6'd36;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,4258,cycle)
    `expect("io_rd_imag",io_rd_imag,-649,cycle)
    `expect("io_rd_real",io_rd_real,4258,cycle)
    `expect("io_rd_imag",io_rd_imag,-649,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd16;
    io_rs1_imag = -39;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,3661,cycle)
    `expect("io_rd_imag",io_rd_imag,-2000,cycle)
    `expect("io_rd_real",io_rd_real,3661,cycle)
    `expect("io_rd_imag",io_rd_imag,-2000,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -10;
    io_rs1_imag = -20;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-273,cycle)
    `expect("io_rd_imag",io_rd_imag,-866,cycle)
    `expect("io_rd_real",io_rd_real,-273,cycle)
    `expect("io_rd_imag",io_rd_imag,-866,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd47;
    io_rs1_imag = 6'd35;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,876,cycle)
    `expect("io_rd_imag",io_rd_imag,-5361,cycle)
    `expect("io_rd_real",io_rd_real,876,cycle)
    `expect("io_rd_imag",io_rd_imag,-5361,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd49;
    io_rs1_imag = -30;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1846,cycle)
    `expect("io_rd_imag",io_rd_imag,-3792,cycle)
    `expect("io_rd_real",io_rd_real,1846,cycle)
    `expect("io_rd_imag",io_rd_imag,-3792,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd40;
    io_rs1_imag = 4'd9;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1928,cycle)
    `expect("io_rd_imag",io_rd_imag,-1689,cycle)
    `expect("io_rd_real",io_rd_real,1928,cycle)
    `expect("io_rd_imag",io_rd_imag,-1689,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = -44;
    io_rs1_imag = -33;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,925,cycle)
    `expect("io_rd_imag",io_rd_imag,-2762,cycle)
    `expect("io_rd_real",io_rd_real,925,cycle)
    `expect("io_rd_imag",io_rd_imag,-2762,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd21;
    io_rs1_imag = -30;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1942,cycle)
    `expect("io_rd_imag",io_rd_imag,-3380,cycle)
    `expect("io_rd_real",io_rd_real,-1942,cycle)
    `expect("io_rd_imag",io_rd_imag,-3380,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd33;
    io_rs1_imag = -34;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-5525,cycle)
    `expect("io_rd_imag",io_rd_imag,-6131,cycle)
    `expect("io_rd_real",io_rd_real,-5525,cycle)
    `expect("io_rd_imag",io_rd_imag,-6131,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 6'd38;
    io_rs1_imag = 3'd6;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1067,cycle)
    `expect("io_rd_imag",io_rd_imag,-4794,cycle)
    `expect("io_rd_real",io_rd_real,1067,cycle)
    `expect("io_rd_imag",io_rd_imag,-4794,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 4'd9;
    io_rs1_imag = -8;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,1019,cycle)
    `expect("io_rd_imag",io_rd_imag,-909,cycle)
    `expect("io_rd_real",io_rd_real,1019,cycle)
    `expect("io_rd_imag",io_rd_imag,-909,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1_real = 5'd20;
    io_rs1_imag = -42;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 7'd91;
    #(1*`CLK_PERIOD)     `expect("io_rd_real",io_rd_real,-1784,cycle)
    `expect("io_rd_imag",io_rd_imag,-2111,cycle)
    `expect("io_rd_real",io_rd_real,-1784,cycle)
    `expect("io_rd_imag",io_rd_imag,-2111,cycle)
    io_valid = 1'd0;

    #`CLK_PERIOD $display("\t **Ran through all test vectors**"); $finish;

  end
endmodule