module SCIEPipelined #(parameter XLEN = 32)(
  input         clock,

  input         valid,
  input  [31:0] insn,
  input  [31:0] rs1,
  input  [31:0] rs2,
  output [31:0] rd
);
reg reset = 0;
  reg [31:0] coeffs_0;
  reg [31:0] coeffs_1;
  reg [31:0] coeffs_2;
  reg [31:0] coeffs_3;
  reg [31:0] coeffs_4;
  reg [31:0] coeffs_5;
  reg [31:0] coeffs_6;
  reg [31:0] coeffs_7;
  reg [31:0] coeffs_8;
  reg [31:0] coeffs_9;
  reg [31:0] coeffs_10;
  reg [31:0] coeffs_11;
  reg [31:0] coeffs_12;
  reg [31:0] coeffs_13;
  reg [31:0] coeffs_14;
  reg [31:0] coeffs_15;
  reg [31:0] coeffs_16;
  reg [31:0] coeffs_17;
  reg [31:0] coeffs_18;
  reg [31:0] coeffs_19;
  reg [31:0] coeffs_20;
  reg [31:0] coeffs_21;
  reg [31:0] coeffs_22;
  reg [31:0] coeffs_23;
  reg [31:0] coeffs_24;
  reg [31:0] coeffs_25;
  reg [31:0] coeffs_26;
  reg [31:0] coeffs_27;
  reg [31:0] coeffs_28;
  reg [31:0] coeffs_29;
  reg [31:0] coeffs_30;
  reg [31:0] coeffs_31;
  reg [31:0] coeffs_32;
  reg [31:0] coeffs_33;
  reg [31:0] coeffs_34;
  reg [31:0] coeffs_35;
  reg [31:0] coeffs_36;
  reg [31:0] coeffs_37;
  reg [31:0] coeffs_38;
  reg [31:0] coeffs_39;
  reg [31:0] coeffs_40;
  reg [31:0] coeffs_41;
  reg [31:0] coeffs_42;
  reg [31:0] coeffs_43;
  reg [31:0] coeffs_44;
  reg [31:0] coeffs_45;
  reg [31:0] coeffs_46;
  reg [31:0] coeffs_47;
  reg [31:0] coeffs_48;
  reg [31:0] coeffs_49;
  reg [31:0] coeffs_50;
  reg [31:0] coeffs_51;
  reg [31:0] coeffs_52;
  reg [31:0] coeffs_53;
  reg [31:0] coeffs_54;
  reg [31:0] coeffs_55;
  reg [31:0] coeffs_56;
  reg [31:0] coeffs_57;
  reg [31:0] coeffs_58;
  reg [31:0] coeffs_59;
  reg [31:0] coeffs_60;
  reg [31:0] coeffs_61;
  reg [31:0] coeffs_62;
  reg [31:0] coeffs_63;
  reg [31:0] coeffs_64;
  reg [31:0] coeffs_65;
  reg [31:0] coeffs_66;
  reg [31:0] coeffs_67;
  reg [31:0] coeffs_68;
  reg [31:0] coeffs_69;
  reg [31:0] coeffs_70;
  reg [31:0] coeffs_71;
  reg [31:0] coeffs_72;
  reg [31:0] coeffs_73;
  reg [31:0] coeffs_74;
  reg [31:0] coeffs_75;
  reg [31:0] coeffs_76;
  reg [31:0] coeffs_77;
  reg [31:0] coeffs_78;
  reg [31:0] coeffs_79;
  reg [31:0] coeffs_80;
  reg [31:0] coeffs_81;
  reg [31:0] coeffs_82;
  reg [31:0] coeffs_83;
  reg [31:0] coeffs_84;
  reg [31:0] coeffs_85;
  reg [31:0] coeffs_86;
  reg [31:0] coeffs_87;
  reg [31:0] coeffs_88;
  reg [31:0] coeffs_89;
  reg [31:0] coeffs_90;
  reg [31:0] coeffs_91;
  reg [31:0] coeffs_92;
  reg [31:0] coeffs_93;
  reg [31:0] coeffs_94;
  reg [31:0] coeffs_95;
  reg [31:0] coeffs_96;
  reg [31:0] coeffs_97;
  reg [31:0] coeffs_98;
  reg [31:0] coeffs_99;
  reg [31:0] coeffs_100;
  reg [31:0] coeffs_101;
  reg [31:0] coeffs_102;
  reg [31:0] coeffs_103;
  reg [31:0] coeffs_104;
  reg [31:0] coeffs_105;
  reg [31:0] coeffs_106;
  reg [31:0] coeffs_107;
  reg [31:0] coeffs_108;
  reg [31:0] coeffs_109;
  reg [31:0] coeffs_110;
  reg [31:0] coeffs_111;
  reg [31:0] coeffs_112;
  reg [31:0] coeffs_113;
  reg [31:0] coeffs_114;
  reg [31:0] coeffs_115;
  reg [31:0] coeffs_116;
  reg [31:0] coeffs_117;
  reg [31:0] coeffs_118;
  reg [31:0] coeffs_119;
  reg [31:0] coeffs_120;
  reg [31:0] coeffs_121;
  reg [31:0] coeffs_122;
  reg [31:0] coeffs_123;
  reg [31:0] coeffs_124;
  reg [31:0] coeffs_125;
  reg [31:0] coeffs_126;
  reg [31:0] coeffs_127;
  reg [31:0] coeffs_128;
  reg [31:0] coeffs_129;
  reg [31:0] coeffs_130;
  reg [31:0] coeffs_131;
  reg [31:0] coeffs_132;
  reg [31:0] coeffs_133;
  reg [31:0] coeffs_134;
  reg [31:0] coeffs_135;
  reg [31:0] coeffs_136;
  reg [31:0] coeffs_137;
  reg [31:0] coeffs_138;
  reg [31:0] coeffs_139;
  reg [31:0] coeffs_140;
  reg [31:0] coeffs_141;
  reg [31:0] coeffs_142;
  reg [31:0] coeffs_143;
  reg [31:0] coeffs_144;
  reg [31:0] coeffs_145;
  reg [31:0] coeffs_146;
  reg [31:0] coeffs_147;
  reg [31:0] coeffs_148;
  reg [31:0] coeffs_149;
  reg [31:0] coeffs_150;
  reg [31:0] coeffs_151;
  reg [31:0] coeffs_152;
  reg [31:0] coeffs_153;
  reg [31:0] coeffs_154;
  reg [31:0] coeffs_155;
  reg [31:0] coeffs_156;
  reg [31:0] coeffs_157;
  reg [31:0] coeffs_158;
  reg [31:0] coeffs_159;
  reg [31:0] coeffs_160;
  reg [31:0] coeffs_161;
  reg [31:0] coeffs_162;
  reg [31:0] coeffs_163;
  reg [31:0] coeffs_164;
  reg [31:0] coeffs_165;
  reg [31:0] coeffs_166;
  reg [31:0] coeffs_167;
  reg [31:0] coeffs_168;
  reg [31:0] coeffs_169;
  reg [31:0] coeffs_170;
  reg [31:0] coeffs_171;
  reg [31:0] coeffs_172;
  reg [31:0] coeffs_173;
  reg [31:0] coeffs_174;
  reg [31:0] coeffs_175;
  reg [31:0] coeffs_176;
  reg [31:0] coeffs_177;
  reg [31:0] coeffs_178;
  reg [31:0] coeffs_179;
  reg [31:0] coeffs_180;
  reg [31:0] coeffs_181;
  reg [31:0] coeffs_182;
  reg [31:0] coeffs_183;
  reg [31:0] coeffs_184;
  reg [31:0] coeffs_185;
  reg [31:0] coeffs_186;
  reg [31:0] coeffs_187;
  reg [31:0] coeffs_188;
  reg [31:0] coeffs_189;
  reg [31:0] coeffs_190;
  reg [31:0] coeffs_191;
  reg [31:0] coeffs_192;
  reg [31:0] coeffs_193;
  reg [31:0] coeffs_194;
  reg [31:0] coeffs_195;
  reg [31:0] coeffs_196;
  reg [31:0] coeffs_197;
  reg [31:0] coeffs_198;
  reg [31:0] coeffs_199;
  reg [31:0] coeffs_200;
  reg [31:0] coeffs_201;
  reg [31:0] coeffs_202;
  reg [31:0] coeffs_203;
  reg [31:0] coeffs_204;
  reg [31:0] coeffs_205;
  reg [31:0] coeffs_206;
  reg [31:0] coeffs_207;
  reg [31:0] coeffs_208;
  reg [31:0] coeffs_209;
  reg [31:0] coeffs_210;
  reg [31:0] coeffs_211;
  reg [31:0] coeffs_212;
  reg [31:0] coeffs_213;
  reg [31:0] coeffs_214;
  reg [31:0] coeffs_215;
  reg [31:0] coeffs_216;
  reg [31:0] coeffs_217;
  reg [31:0] coeffs_218;
  reg [31:0] coeffs_219;
  reg [31:0] coeffs_220;
  reg [31:0] coeffs_221;
  reg [31:0] coeffs_222;
  reg [31:0] coeffs_223;
  reg [31:0] coeffs_224;
  reg [31:0] coeffs_225;
  reg [31:0] coeffs_226;
  reg [31:0] coeffs_227;
  reg [31:0] coeffs_228;
  reg [31:0] coeffs_229;
  reg [31:0] coeffs_230;
  reg [31:0] coeffs_231;
  reg [31:0] coeffs_232;
  reg [31:0] coeffs_233;
  reg [31:0] coeffs_234;
  reg [31:0] coeffs_235;
  reg [31:0] coeffs_236;
  reg [31:0] coeffs_237;
  reg [31:0] coeffs_238;
  reg [31:0] coeffs_239;
  reg [31:0] coeffs_240;
  reg [31:0] coeffs_241;
  reg [31:0] coeffs_242;
  reg [31:0] coeffs_243;
  reg [31:0] coeffs_244;
  reg [31:0] coeffs_245;
  reg [31:0] coeffs_246;
  reg [31:0] coeffs_247;
  reg [31:0] coeffs_248;
  reg [31:0] coeffs_249;
  reg [31:0] coeffs_250;
  reg [31:0] coeffs_251;
  reg [31:0] coeffs_252;
  reg [31:0] coeffs_253;
  reg [31:0] coeffs_254;
  reg [31:0] coeffs_255;
  reg [31:0] coeffs_256;
  reg [31:0] coeffs_257;
  reg [31:0] coeffs_258;
  reg [31:0] coeffs_259;
  reg [31:0] coeffs_260;
  reg [31:0] coeffs_261;
  reg [31:0] coeffs_262;
  reg [31:0] coeffs_263;
  reg [31:0] coeffs_264;
  reg [31:0] coeffs_265;
  reg [31:0] coeffs_266;
  reg [31:0] coeffs_267;
  reg [31:0] coeffs_268;
  reg [31:0] coeffs_269;
  reg [31:0] coeffs_270;
  reg [31:0] coeffs_271;
  reg [31:0] coeffs_272;
  reg [31:0] coeffs_273;
  reg [31:0] coeffs_274;
  reg [31:0] coeffs_275;
  reg [31:0] coeffs_276;
  reg [31:0] coeffs_277;
  reg [31:0] coeffs_278;
  reg [31:0] coeffs_279;
  reg [31:0] coeffs_280;
  reg [31:0] coeffs_281;
  reg [31:0] coeffs_282;
  reg [31:0] coeffs_283;
  reg [31:0] coeffs_284;
  reg [31:0] coeffs_285;
  reg [31:0] coeffs_286;
  reg [31:0] coeffs_287;
  reg [31:0] coeffs_288;
  reg [31:0] coeffs_289;
  reg [31:0] coeffs_290;
  reg [31:0] coeffs_291;
  reg [31:0] coeffs_292;
  reg [31:0] coeffs_293;
  reg [31:0] coeffs_294;
  reg [31:0] coeffs_295;
  reg [31:0] coeffs_296;
  reg [31:0] coeffs_297;
  reg [31:0] coeffs_298;
  reg [31:0] coeffs_299;
  reg [31:0] coeffs_300;
  reg [31:0] coeffs_301;
  reg [31:0] coeffs_302;
  reg [31:0] coeffs_303;
  reg [31:0] coeffs_304;
  reg [31:0] coeffs_305;
  reg [31:0] coeffs_306;
  reg [31:0] coeffs_307;
  reg [31:0] coeffs_308;
  reg [31:0] coeffs_309;
  reg [31:0] coeffs_310;
  reg [31:0] coeffs_311;
  reg [31:0] coeffs_312;
  reg [31:0] coeffs_313;
  reg [31:0] coeffs_314;
  reg [31:0] coeffs_315;
  reg [31:0] coeffs_316;
  reg [31:0] coeffs_317;
  reg [31:0] coeffs_318;
  reg [31:0] coeffs_319;
  reg [31:0] coeffs_320;
  reg [31:0] coeffs_321;
  reg [31:0] coeffs_322;
  reg [31:0] coeffs_323;
  reg [31:0] coeffs_324;
  reg [31:0] coeffs_325;
  reg [31:0] coeffs_326;
  reg [31:0] coeffs_327;
  reg [31:0] coeffs_328;
  reg [31:0] coeffs_329;
  reg [31:0] coeffs_330;
  reg [31:0] coeffs_331;
  reg [31:0] coeffs_332;
  reg [31:0] coeffs_333;
  reg [31:0] coeffs_334;
  reg [31:0] coeffs_335;
  reg [31:0] coeffs_336;
  reg [31:0] coeffs_337;
  reg [31:0] coeffs_338;
  reg [31:0] coeffs_339;
  reg [31:0] coeffs_340;
  reg [31:0] coeffs_341;
  reg [31:0] coeffs_342;
  reg [31:0] coeffs_343;
  reg [31:0] coeffs_344;
  reg [31:0] coeffs_345;
  reg [31:0] coeffs_346;
  reg [31:0] coeffs_347;
  reg [31:0] coeffs_348;
  reg [31:0] coeffs_349;
  reg [31:0] coeffs_350;
  reg [31:0] coeffs_351;
  reg [31:0] coeffs_352;
  reg [31:0] coeffs_353;
  reg [31:0] coeffs_354;
  reg [31:0] coeffs_355;
  reg [31:0] coeffs_356;
  reg [31:0] coeffs_357;
  reg [31:0] coeffs_358;
  reg [31:0] coeffs_359;
  reg [31:0] coeffs_360;
  reg [31:0] coeffs_361;
  reg [31:0] coeffs_362;
  reg [31:0] coeffs_363;
  reg [31:0] coeffs_364;
  reg [31:0] coeffs_365;
  reg [31:0] coeffs_366;
  reg [31:0] coeffs_367;
  reg [31:0] coeffs_368;
  reg [31:0] coeffs_369;
  reg [31:0] coeffs_370;
  reg [31:0] coeffs_371;
  reg [31:0] coeffs_372;
  reg [31:0] coeffs_373;
  reg [31:0] coeffs_374;
  reg [31:0] coeffs_375;
  reg [31:0] coeffs_376;
  reg [31:0] coeffs_377;
  reg [31:0] coeffs_378;
  reg [31:0] coeffs_379;
  reg [31:0] coeffs_380;
  reg [31:0] coeffs_381;
  reg [31:0] coeffs_382;
  reg [31:0] coeffs_383;
  reg [31:0] coeffs_384;
  reg [31:0] coeffs_385;
  reg [31:0] coeffs_386;
  reg [31:0] coeffs_387;
  reg [31:0] coeffs_388;
  reg [31:0] coeffs_389;
  reg [31:0] coeffs_390;
  reg [31:0] coeffs_391;
  reg [31:0] coeffs_392;
  reg [31:0] coeffs_393;
  reg [31:0] coeffs_394;
  reg [31:0] coeffs_395;
  reg [31:0] coeffs_396;
  reg [31:0] coeffs_397;
  reg [31:0] coeffs_398;
  reg [31:0] coeffs_399;
  reg [31:0] coeffs_400;
  reg [31:0] coeffs_401;
  reg [31:0] coeffs_402;
  reg [31:0] coeffs_403;
  reg [31:0] coeffs_404;
  reg [31:0] coeffs_405;
  reg [31:0] coeffs_406;
  reg [31:0] coeffs_407;
  reg [31:0] coeffs_408;
  reg [31:0] coeffs_409;
  reg [31:0] coeffs_410;
  reg [31:0] coeffs_411;
  reg [31:0] coeffs_412;
  reg [31:0] coeffs_413;
  reg [31:0] coeffs_414;
  reg [31:0] coeffs_415;
  reg [31:0] coeffs_416;
  reg [31:0] coeffs_417;
  reg [31:0] coeffs_418;
  reg [31:0] coeffs_419;
  reg [31:0] coeffs_420;
  reg [31:0] coeffs_421;
  reg [31:0] coeffs_422;
  reg [31:0] coeffs_423;
  reg [31:0] coeffs_424;
  reg [31:0] coeffs_425;
  reg [31:0] coeffs_426;
  reg [31:0] coeffs_427;
  reg [31:0] coeffs_428;
  reg [31:0] coeffs_429;
  reg [31:0] coeffs_430;
  reg [31:0] coeffs_431;
  reg [31:0] coeffs_432;
  reg [31:0] coeffs_433;
  reg [31:0] coeffs_434;
  reg [31:0] coeffs_435;
  reg [31:0] coeffs_436;
  reg [31:0] coeffs_437;
  reg [31:0] coeffs_438;
  reg [31:0] coeffs_439;
  reg [31:0] coeffs_440;
  reg [31:0] coeffs_441;
  reg [31:0] coeffs_442;
  reg [31:0] coeffs_443;
  reg [31:0] coeffs_444;
  reg [31:0] coeffs_445;
  reg [31:0] coeffs_446;
  reg [31:0] coeffs_447;
  reg [31:0] coeffs_448;
  reg [31:0] coeffs_449;
  reg [31:0] coeffs_450;
  reg [31:0] coeffs_451;
  reg [31:0] coeffs_452;
  reg [31:0] coeffs_453;
  reg [31:0] coeffs_454;
  reg [31:0] coeffs_455;
  reg [31:0] coeffs_456;
  reg [31:0] coeffs_457;
  reg [31:0] coeffs_458;
  reg [31:0] coeffs_459;
  reg [31:0] coeffs_460;
  reg [31:0] coeffs_461;
  reg [31:0] coeffs_462;
  reg [31:0] coeffs_463;
  reg [31:0] coeffs_464;
  reg [31:0] coeffs_465;
  reg [31:0] coeffs_466;
  reg [31:0] coeffs_467;
  reg [31:0] coeffs_468;
  reg [31:0] coeffs_469;
  reg [31:0] coeffs_470;
  reg [31:0] coeffs_471;
  reg [31:0] coeffs_472;
  reg [31:0] coeffs_473;
  reg [31:0] coeffs_474;
  reg [31:0] coeffs_475;
  reg [31:0] coeffs_476;
  reg [31:0] coeffs_477;
  reg [31:0] coeffs_478;
  reg [31:0] coeffs_479;
  reg [31:0] coeffs_480;
  reg [31:0] coeffs_481;
  reg [31:0] coeffs_482;
  reg [31:0] coeffs_483;
  reg [31:0] coeffs_484;
  reg [31:0] coeffs_485;
  reg [31:0] coeffs_486;
  reg [31:0] coeffs_487;
  reg [31:0] coeffs_488;
  reg [31:0] coeffs_489;
  reg [31:0] coeffs_490;
  reg [31:0] coeffs_491;
  reg [31:0] coeffs_492;
  reg [31:0] coeffs_493;
  reg [31:0] coeffs_494;
  reg [31:0] coeffs_495;
  reg [31:0] coeffs_496;
  reg [31:0] coeffs_497;
  reg [31:0] coeffs_498;
  reg [31:0] coeffs_499;
  reg [31:0] coeffs_500;
  reg [31:0] coeffs_501;
  reg [31:0] coeffs_502;
  reg [31:0] coeffs_503;
  reg [31:0] coeffs_504;
  reg [31:0] coeffs_505;
  reg [31:0] coeffs_506;
  reg [31:0] coeffs_507;
  reg [31:0] coeffs_508;
  reg [31:0] coeffs_509;
  reg [31:0] coeffs_510;
  reg [31:0] coeffs_511;
  reg [31:0] coeffs_512;
  reg [31:0] coeffs_513;
  reg [31:0] coeffs_514;
  reg [31:0] coeffs_515;
  reg [31:0] coeffs_516;
  reg [31:0] coeffs_517;
  reg [31:0] coeffs_518;
  reg [31:0] coeffs_519;
  reg [31:0] coeffs_520;
  reg [31:0] coeffs_521;
  reg [31:0] coeffs_522;
  reg [31:0] coeffs_523;
  reg [31:0] coeffs_524;
  reg [31:0] coeffs_525;
  reg [31:0] coeffs_526;
  reg [31:0] coeffs_527;
  reg [31:0] coeffs_528;
  reg [31:0] coeffs_529;
  reg [31:0] coeffs_530;
  reg [31:0] coeffs_531;
  reg [31:0] coeffs_532;
  reg [31:0] coeffs_533;
  reg [31:0] coeffs_534;
  reg [31:0] coeffs_535;
  reg [31:0] coeffs_536;
  reg [31:0] coeffs_537;
  reg [31:0] coeffs_538;
  reg [31:0] coeffs_539;
  reg [31:0] coeffs_540;
  reg [31:0] coeffs_541;
  reg [31:0] coeffs_542;
  reg [31:0] coeffs_543;
  reg [31:0] coeffs_544;
  reg [31:0] coeffs_545;
  reg [31:0] coeffs_546;
  reg [31:0] coeffs_547;
  reg [31:0] coeffs_548;
  reg [31:0] coeffs_549;
  reg [31:0] coeffs_550;
  reg [31:0] coeffs_551;
  reg [31:0] coeffs_552;
  reg [31:0] coeffs_553;
  reg [31:0] coeffs_554;
  reg [31:0] coeffs_555;
  reg [31:0] coeffs_556;
  reg [31:0] coeffs_557;
  reg [31:0] coeffs_558;
  reg [31:0] coeffs_559;
  reg [31:0] coeffs_560;
  reg [31:0] coeffs_561;
  reg [31:0] coeffs_562;
  reg [31:0] coeffs_563;
  reg [31:0] coeffs_564;
  reg [31:0] coeffs_565;
  reg [31:0] coeffs_566;
  reg [31:0] coeffs_567;
  reg [31:0] coeffs_568;
  reg [31:0] coeffs_569;
  reg [31:0] coeffs_570;
  reg [31:0] coeffs_571;
  reg [31:0] coeffs_572;
  reg [31:0] coeffs_573;
  reg [31:0] coeffs_574;
  reg [31:0] coeffs_575;
  reg [31:0] coeffs_576;
  reg [31:0] coeffs_577;
  reg [31:0] coeffs_578;
  reg [31:0] coeffs_579;
  reg [31:0] coeffs_580;
  reg [31:0] coeffs_581;
  reg [31:0] coeffs_582;
  reg [31:0] coeffs_583;
  reg [31:0] coeffs_584;
  reg [31:0] coeffs_585;
  reg [31:0] coeffs_586;
  reg [31:0] coeffs_587;
  reg [31:0] coeffs_588;
  reg [31:0] coeffs_589;
  reg [31:0] coeffs_590;
  reg [31:0] coeffs_591;
  reg [31:0] coeffs_592;
  reg [31:0] coeffs_593;
  reg [31:0] coeffs_594;
  reg [31:0] coeffs_595;
  reg [31:0] coeffs_596;
  reg [31:0] coeffs_597;
  reg [31:0] coeffs_598;
  reg [31:0] coeffs_599;
  reg [31:0] coeffs_600;
  reg [31:0] coeffs_601;
  reg [31:0] coeffs_602;
  reg [31:0] coeffs_603;
  reg [31:0] coeffs_604;
  reg [31:0] coeffs_605;
  reg [31:0] coeffs_606;
  reg [31:0] coeffs_607;
  reg [31:0] coeffs_608;
  reg [31:0] coeffs_609;
  reg [31:0] coeffs_610;
  reg [31:0] coeffs_611;
  reg [31:0] coeffs_612;
  reg [31:0] coeffs_613;
  reg [31:0] coeffs_614;
  reg [31:0] coeffs_615;
  reg [31:0] coeffs_616;
  reg [31:0] coeffs_617;
  reg [31:0] coeffs_618;
  reg [31:0] coeffs_619;
  reg [31:0] coeffs_620;
  reg [31:0] coeffs_621;
  reg [31:0] coeffs_622;
  reg [31:0] coeffs_623;
  reg [31:0] coeffs_624;
  reg [31:0] coeffs_625;
  reg [31:0] coeffs_626;
  reg [31:0] coeffs_627;
  reg [31:0] coeffs_628;
  reg [31:0] coeffs_629;
  reg [31:0] coeffs_630;
  reg [31:0] coeffs_631;
  reg [31:0] coeffs_632;
  reg [31:0] coeffs_633;
  reg [31:0] coeffs_634;
  reg [31:0] coeffs_635;
  reg [31:0] coeffs_636;
  reg [31:0] coeffs_637;
  reg [31:0] coeffs_638;
  reg [31:0] coeffs_639;
  reg [31:0] coeffs_640;
  reg [31:0] coeffs_641;
  reg [31:0] coeffs_642;
  reg [31:0] coeffs_643;
  reg [31:0] coeffs_644;
  reg [31:0] coeffs_645;
  reg [31:0] coeffs_646;
  reg [31:0] coeffs_647;
  reg [31:0] coeffs_648;
  reg [31:0] coeffs_649;
  reg [31:0] coeffs_650;
  reg [31:0] coeffs_651;
  reg [31:0] coeffs_652;
  reg [31:0] coeffs_653;
  reg [31:0] coeffs_654;
  reg [31:0] coeffs_655;
  reg [31:0] coeffs_656;
  reg [31:0] coeffs_657;
  reg [31:0] coeffs_658;
  reg [31:0] coeffs_659;
  reg [31:0] coeffs_660;
  reg [31:0] coeffs_661;
  reg [31:0] coeffs_662;
  reg [31:0] coeffs_663;
  reg [31:0] coeffs_664;
  reg [31:0] coeffs_665;
  reg [31:0] coeffs_666;
  reg [31:0] coeffs_667;
  reg [31:0] coeffs_668;
  reg [31:0] coeffs_669;
  reg [31:0] coeffs_670;
  reg [31:0] coeffs_671;
  reg [31:0] coeffs_672;
  reg [31:0] coeffs_673;
  reg [31:0] coeffs_674;
  reg [31:0] coeffs_675;
  reg [31:0] coeffs_676;
  reg [31:0] coeffs_677;
  reg [31:0] coeffs_678;
  reg [31:0] coeffs_679;
  reg [31:0] coeffs_680;
  reg [31:0] coeffs_681;
  reg [31:0] coeffs_682;
  reg [31:0] coeffs_683;
  reg [31:0] coeffs_684;
  reg [31:0] coeffs_685;
  reg [31:0] coeffs_686;
  reg [31:0] coeffs_687;
  reg [31:0] coeffs_688;
  reg [31:0] coeffs_689;
  reg [31:0] coeffs_690;
  reg [31:0] coeffs_691;
  reg [31:0] coeffs_692;
  reg [31:0] coeffs_693;
  reg [31:0] coeffs_694;
  reg [31:0] coeffs_695;
  reg [31:0] coeffs_696;
  reg [31:0] coeffs_697;
  reg [31:0] coeffs_698;
  reg [31:0] coeffs_699;
  reg [31:0] coeffs_700;
  reg [31:0] coeffs_701;
  reg [31:0] coeffs_702;
  reg [31:0] coeffs_703;
  reg [31:0] coeffs_704;
  reg [31:0] coeffs_705;
  reg [31:0] coeffs_706;
  reg [31:0] coeffs_707;
  reg [31:0] coeffs_708;
  reg [31:0] coeffs_709;
  reg [31:0] coeffs_710;
  reg [31:0] coeffs_711;
  reg [31:0] coeffs_712;
  reg [31:0] coeffs_713;
  reg [31:0] coeffs_714;
  reg [31:0] coeffs_715;
  reg [31:0] coeffs_716;
  reg [31:0] coeffs_717;
  reg [31:0] coeffs_718;
  reg [31:0] coeffs_719;
  reg [31:0] coeffs_720;
  reg [31:0] coeffs_721;
  reg [31:0] coeffs_722;
  reg [31:0] coeffs_723;
  reg [31:0] coeffs_724;
  reg [31:0] coeffs_725;
  reg [31:0] coeffs_726;
  reg [31:0] coeffs_727;
  reg [31:0] coeffs_728;
  reg [31:0] coeffs_729;
  reg [31:0] coeffs_730;
  reg [31:0] coeffs_731;
  reg [31:0] coeffs_732;
  reg [31:0] coeffs_733;
  reg [31:0] coeffs_734;
  reg [31:0] coeffs_735;
  reg [31:0] coeffs_736;
  reg [31:0] coeffs_737;
  reg [31:0] coeffs_738;
  reg [31:0] coeffs_739;
  reg [31:0] coeffs_740;
  reg [31:0] coeffs_741;
  reg [31:0] coeffs_742;
  reg [31:0] coeffs_743;
  reg [31:0] coeffs_744;
  reg [31:0] coeffs_745;
  reg [31:0] coeffs_746;
  reg [31:0] coeffs_747;
  reg [31:0] coeffs_748;
  reg [31:0] coeffs_749;
  reg [31:0] coeffs_750;
  reg [31:0] coeffs_751;
  reg [31:0] coeffs_752;
  reg [31:0] coeffs_753;
  reg [31:0] coeffs_754;
  reg [31:0] coeffs_755;
  reg [31:0] coeffs_756;
  reg [31:0] coeffs_757;
  reg [31:0] coeffs_758;
  reg [31:0] coeffs_759;
  reg [31:0] coeffs_760;
  reg [31:0] coeffs_761;
  reg [31:0] coeffs_762;
  reg [31:0] coeffs_763;
  reg [31:0] coeffs_764;
  reg [31:0] coeffs_765;
  reg [31:0] coeffs_766;
  reg [31:0] coeffs_767;
  reg [31:0] coeffs_768;
  reg [31:0] coeffs_769;
  reg [31:0] coeffs_770;
  reg [31:0] coeffs_771;
  reg [31:0] coeffs_772;
  reg [31:0] coeffs_773;
  reg [31:0] coeffs_774;
  reg [31:0] coeffs_775;
  reg [31:0] coeffs_776;
  reg [31:0] coeffs_777;
  reg [31:0] coeffs_778;
  reg [31:0] coeffs_779;
  reg [31:0] coeffs_780;
  reg [31:0] coeffs_781;
  reg [31:0] coeffs_782;
  reg [31:0] coeffs_783;
  reg [31:0] coeffs_784;
  reg [31:0] coeffs_785;
  reg [31:0] coeffs_786;
  reg [31:0] coeffs_787;
  reg [31:0] coeffs_788;
  reg [31:0] coeffs_789;
  reg [31:0] coeffs_790;
  reg [31:0] coeffs_791;
  reg [31:0] coeffs_792;
  reg [31:0] coeffs_793;
  reg [31:0] coeffs_794;
  reg [31:0] coeffs_795;
  reg [31:0] coeffs_796;
  reg [31:0] coeffs_797;
  reg [31:0] coeffs_798;
  reg [31:0] coeffs_799;
  reg [31:0] coeffs_800;
  reg [31:0] coeffs_801;
  reg [31:0] coeffs_802;
  reg [31:0] coeffs_803;
  reg [31:0] coeffs_804;
  reg [31:0] coeffs_805;
  reg [31:0] coeffs_806;
  reg [31:0] coeffs_807;
  reg [31:0] coeffs_808;
  reg [31:0] coeffs_809;
  reg [31:0] coeffs_810;
  reg [31:0] coeffs_811;
  reg [31:0] coeffs_812;
  reg [31:0] coeffs_813;
  reg [31:0] coeffs_814;
  reg [31:0] coeffs_815;
  reg [31:0] coeffs_816;
  reg [31:0] coeffs_817;
  reg [31:0] coeffs_818;
  reg [31:0] coeffs_819;
  reg [31:0] coeffs_820;
  reg [31:0] coeffs_821;
  reg [31:0] coeffs_822;
  reg [31:0] coeffs_823;
  reg [31:0] coeffs_824;
  reg [31:0] coeffs_825;
  reg [31:0] coeffs_826;
  reg [31:0] coeffs_827;
  reg [31:0] coeffs_828;
  reg [31:0] coeffs_829;
  reg [31:0] coeffs_830;
  reg [31:0] coeffs_831;
  reg [31:0] coeffs_832;
  reg [31:0] coeffs_833;
  reg [31:0] coeffs_834;
  reg [31:0] coeffs_835;
  reg [31:0] coeffs_836;
  reg [31:0] coeffs_837;
  reg [31:0] coeffs_838;
  reg [31:0] coeffs_839;
  reg [31:0] coeffs_840;
  reg [31:0] coeffs_841;
  reg [31:0] coeffs_842;
  reg [31:0] coeffs_843;
  reg [31:0] coeffs_844;
  reg [31:0] coeffs_845;
  reg [31:0] coeffs_846;
  reg [31:0] coeffs_847;
  reg [31:0] coeffs_848;
  reg [31:0] coeffs_849;
  reg [31:0] coeffs_850;
  reg [31:0] coeffs_851;
  reg [31:0] coeffs_852;
  reg [31:0] coeffs_853;
  reg [31:0] coeffs_854;
  reg [31:0] coeffs_855;
  reg [31:0] coeffs_856;
  reg [31:0] coeffs_857;
  reg [31:0] coeffs_858;
  reg [31:0] coeffs_859;
  reg [31:0] coeffs_860;
  reg [31:0] coeffs_861;
  reg [31:0] coeffs_862;
  reg [31:0] coeffs_863;
  reg [31:0] coeffs_864;
  reg [31:0] coeffs_865;
  reg [31:0] coeffs_866;
  reg [31:0] coeffs_867;
  reg [31:0] coeffs_868;
  reg [31:0] coeffs_869;
  reg [31:0] coeffs_870;
  reg [31:0] coeffs_871;
  reg [31:0] coeffs_872;
  reg [31:0] coeffs_873;
  reg [31:0] coeffs_874;
  reg [31:0] coeffs_875;
  reg [31:0] coeffs_876;
  reg [31:0] coeffs_877;
  reg [31:0] coeffs_878;
  reg [31:0] coeffs_879;
  reg [31:0] coeffs_880;
  reg [31:0] coeffs_881;
  reg [31:0] coeffs_882;
  reg [31:0] coeffs_883;
  reg [31:0] coeffs_884;
  reg [31:0] coeffs_885;
  reg [31:0] coeffs_886;
  reg [31:0] coeffs_887;
  reg [31:0] coeffs_888;
  reg [31:0] coeffs_889;
  reg [31:0] coeffs_890;
  reg [31:0] coeffs_891;
  reg [31:0] coeffs_892;
  reg [31:0] coeffs_893;
  reg [31:0] coeffs_894;
  reg [31:0] coeffs_895;
  reg [31:0] coeffs_896;
  reg [31:0] coeffs_897;
  reg [31:0] coeffs_898;
  reg [31:0] coeffs_899;
  reg [31:0] coeffs_900;
  reg [31:0] coeffs_901;
  reg [31:0] coeffs_902;
  reg [31:0] coeffs_903;
  reg [31:0] coeffs_904;
  reg [31:0] coeffs_905;
  reg [31:0] coeffs_906;
  reg [31:0] coeffs_907;
  reg [31:0] coeffs_908;
  reg [31:0] coeffs_909;
  reg [31:0] coeffs_910;
  reg [31:0] coeffs_911;
  reg [31:0] coeffs_912;
  reg [31:0] coeffs_913;
  reg [31:0] coeffs_914;
  reg [31:0] coeffs_915;
  reg [31:0] coeffs_916;
  reg [31:0] coeffs_917;
  reg [31:0] coeffs_918;
  reg [31:0] coeffs_919;
  reg [31:0] coeffs_920;
  reg [31:0] coeffs_921;
  reg [31:0] coeffs_922;
  reg [31:0] coeffs_923;
  reg [31:0] coeffs_924;
  reg [31:0] coeffs_925;
  reg [31:0] coeffs_926;
  reg [31:0] coeffs_927;
  reg [31:0] coeffs_928;
  reg [31:0] coeffs_929;
  reg [31:0] coeffs_930;
  reg [31:0] coeffs_931;
  reg [31:0] coeffs_932;
  reg [31:0] coeffs_933;
  reg [31:0] coeffs_934;
  reg [31:0] coeffs_935;
  reg [31:0] coeffs_936;
  reg [31:0] coeffs_937;
  reg [31:0] coeffs_938;
  reg [31:0] coeffs_939;
  reg [31:0] coeffs_940;
  reg [31:0] coeffs_941;
  reg [31:0] coeffs_942;
  reg [31:0] coeffs_943;
  reg [31:0] coeffs_944;
  reg [31:0] coeffs_945;
  reg [31:0] coeffs_946;
  reg [31:0] coeffs_947;
  reg [31:0] coeffs_948;
  reg [31:0] coeffs_949;
  reg [31:0] coeffs_950;
  reg [31:0] coeffs_951;
  reg [31:0] coeffs_952;
  reg [31:0] coeffs_953;
  reg [31:0] coeffs_954;
  reg [31:0] coeffs_955;
  reg [31:0] coeffs_956;
  reg [31:0] coeffs_957;
  reg [31:0] coeffs_958;
  reg [31:0] coeffs_959;
  reg [31:0] coeffs_960;
  reg [31:0] coeffs_961;
  reg [31:0] coeffs_962;
  reg [31:0] coeffs_963;
  reg [31:0] coeffs_964;
  reg [31:0] coeffs_965;
  reg [31:0] coeffs_966;
  reg [31:0] coeffs_967;
  reg [31:0] coeffs_968;
  reg [31:0] coeffs_969;
  reg [31:0] coeffs_970;
  reg [31:0] coeffs_971;
  reg [31:0] coeffs_972;
  reg [31:0] coeffs_973;
  reg [31:0] coeffs_974;
  reg [31:0] coeffs_975;
  reg [31:0] coeffs_976;
  reg [31:0] coeffs_977;
  reg [31:0] coeffs_978;
  reg [31:0] coeffs_979;
  reg [31:0] coeffs_980;
  reg [31:0] coeffs_981;
  reg [31:0] coeffs_982;
  reg [31:0] coeffs_983;
  reg [31:0] coeffs_984;
  reg [31:0] coeffs_985;
  reg [31:0] coeffs_986;
  reg [31:0] coeffs_987;
  reg [31:0] coeffs_988;
  reg [31:0] coeffs_989;
  reg [31:0] coeffs_990;
  reg [31:0] coeffs_991;
  reg [31:0] coeffs_992;
  reg [31:0] coeffs_993;
  reg [31:0] coeffs_994;
  reg [31:0] coeffs_995;
  reg [31:0] coeffs_996;
  reg [31:0] coeffs_997;
  reg [31:0] coeffs_998;
  reg [31:0] coeffs_999;
  reg [31:0] data_0;
  reg [31:0] data_1;
  reg [31:0] data_2;
  reg [31:0] data_3;
  reg [31:0] data_4;
  reg [31:0] data_5;
  reg [31:0] data_6;
  reg [31:0] data_7;
  reg [31:0] data_8;
  reg [31:0] data_9;
  reg [31:0] data_10;
  reg [31:0] data_11;
  reg [31:0] data_12;
  reg [31:0] data_13;
  reg [31:0] data_14;
  reg [31:0] data_15;
  reg [31:0] data_16;
  reg [31:0] data_17;
  reg [31:0] data_18;
  reg [31:0] data_19;
  reg [31:0] data_20;
  reg [31:0] data_21;
  reg [31:0] data_22;
  reg [31:0] data_23;
  reg [31:0] data_24;
  reg [31:0] data_25;
  reg [31:0] data_26;
  reg [31:0] data_27;
  reg [31:0] data_28;
  reg [31:0] data_29;
  reg [31:0] data_30;
  reg [31:0] data_31;
  reg [31:0] data_32;
  reg [31:0] data_33;
  reg [31:0] data_34;
  reg [31:0] data_35;
  reg [31:0] data_36;
  reg [31:0] data_37;
  reg [31:0] data_38;
  reg [31:0] data_39;
  reg [31:0] data_40;
  reg [31:0] data_41;
  reg [31:0] data_42;
  reg [31:0] data_43;
  reg [31:0] data_44;
  reg [31:0] data_45;
  reg [31:0] data_46;
  reg [31:0] data_47;
  reg [31:0] data_48;
  reg [31:0] data_49;
  reg [31:0] data_50;
  reg [31:0] data_51;
  reg [31:0] data_52;
  reg [31:0] data_53;
  reg [31:0] data_54;
  reg [31:0] data_55;
  reg [31:0] data_56;
  reg [31:0] data_57;
  reg [31:0] data_58;
  reg [31:0] data_59;
  reg [31:0] data_60;
  reg [31:0] data_61;
  reg [31:0] data_62;
  reg [31:0] data_63;
  reg [31:0] data_64;
  reg [31:0] data_65;
  reg [31:0] data_66;
  reg [31:0] data_67;
  reg [31:0] data_68;
  reg [31:0] data_69;
  reg [31:0] data_70;
  reg [31:0] data_71;
  reg [31:0] data_72;
  reg [31:0] data_73;
  reg [31:0] data_74;
  reg [31:0] data_75;
  reg [31:0] data_76;
  reg [31:0] data_77;
  reg [31:0] data_78;
  reg [31:0] data_79;
  reg [31:0] data_80;
  reg [31:0] data_81;
  reg [31:0] data_82;
  reg [31:0] data_83;
  reg [31:0] data_84;
  reg [31:0] data_85;
  reg [31:0] data_86;
  reg [31:0] data_87;
  reg [31:0] data_88;
  reg [31:0] data_89;
  reg [31:0] data_90;
  reg [31:0] data_91;
  reg [31:0] data_92;
  reg [31:0] data_93;
  reg [31:0] data_94;
  reg [31:0] data_95;
  reg [31:0] data_96;
  reg [31:0] data_97;
  reg [31:0] data_98;
  reg [31:0] data_99;
  reg [31:0] data_100;
  reg [31:0] data_101;
  reg [31:0] data_102;
  reg [31:0] data_103;
  reg [31:0] data_104;
  reg [31:0] data_105;
  reg [31:0] data_106;
  reg [31:0] data_107;
  reg [31:0] data_108;
  reg [31:0] data_109;
  reg [31:0] data_110;
  reg [31:0] data_111;
  reg [31:0] data_112;
  reg [31:0] data_113;
  reg [31:0] data_114;
  reg [31:0] data_115;
  reg [31:0] data_116;
  reg [31:0] data_117;
  reg [31:0] data_118;
  reg [31:0] data_119;
  reg [31:0] data_120;
  reg [31:0] data_121;
  reg [31:0] data_122;
  reg [31:0] data_123;
  reg [31:0] data_124;
  reg [31:0] data_125;
  reg [31:0] data_126;
  reg [31:0] data_127;
  reg [31:0] data_128;
  reg [31:0] data_129;
  reg [31:0] data_130;
  reg [31:0] data_131;
  reg [31:0] data_132;
  reg [31:0] data_133;
  reg [31:0] data_134;
  reg [31:0] data_135;
  reg [31:0] data_136;
  reg [31:0] data_137;
  reg [31:0] data_138;
  reg [31:0] data_139;
  reg [31:0] data_140;
  reg [31:0] data_141;
  reg [31:0] data_142;
  reg [31:0] data_143;
  reg [31:0] data_144;
  reg [31:0] data_145;
  reg [31:0] data_146;
  reg [31:0] data_147;
  reg [31:0] data_148;
  reg [31:0] data_149;
  reg [31:0] data_150;
  reg [31:0] data_151;
  reg [31:0] data_152;
  reg [31:0] data_153;
  reg [31:0] data_154;
  reg [31:0] data_155;
  reg [31:0] data_156;
  reg [31:0] data_157;
  reg [31:0] data_158;
  reg [31:0] data_159;
  reg [31:0] data_160;
  reg [31:0] data_161;
  reg [31:0] data_162;
  reg [31:0] data_163;
  reg [31:0] data_164;
  reg [31:0] data_165;
  reg [31:0] data_166;
  reg [31:0] data_167;
  reg [31:0] data_168;
  reg [31:0] data_169;
  reg [31:0] data_170;
  reg [31:0] data_171;
  reg [31:0] data_172;
  reg [31:0] data_173;
  reg [31:0] data_174;
  reg [31:0] data_175;
  reg [31:0] data_176;
  reg [31:0] data_177;
  reg [31:0] data_178;
  reg [31:0] data_179;
  reg [31:0] data_180;
  reg [31:0] data_181;
  reg [31:0] data_182;
  reg [31:0] data_183;
  reg [31:0] data_184;
  reg [31:0] data_185;
  reg [31:0] data_186;
  reg [31:0] data_187;
  reg [31:0] data_188;
  reg [31:0] data_189;
  reg [31:0] data_190;
  reg [31:0] data_191;
  reg [31:0] data_192;
  reg [31:0] data_193;
  reg [31:0] data_194;
  reg [31:0] data_195;
  reg [31:0] data_196;
  reg [31:0] data_197;
  reg [31:0] data_198;
  reg [31:0] data_199;
  reg [31:0] data_200;
  reg [31:0] data_201;
  reg [31:0] data_202;
  reg [31:0] data_203;
  reg [31:0] data_204;
  reg [31:0] data_205;
  reg [31:0] data_206;
  reg [31:0] data_207;
  reg [31:0] data_208;
  reg [31:0] data_209;
  reg [31:0] data_210;
  reg [31:0] data_211;
  reg [31:0] data_212;
  reg [31:0] data_213;
  reg [31:0] data_214;
  reg [31:0] data_215;
  reg [31:0] data_216;
  reg [31:0] data_217;
  reg [31:0] data_218;
  reg [31:0] data_219;
  reg [31:0] data_220;
  reg [31:0] data_221;
  reg [31:0] data_222;
  reg [31:0] data_223;
  reg [31:0] data_224;
  reg [31:0] data_225;
  reg [31:0] data_226;
  reg [31:0] data_227;
  reg [31:0] data_228;
  reg [31:0] data_229;
  reg [31:0] data_230;
  reg [31:0] data_231;
  reg [31:0] data_232;
  reg [31:0] data_233;
  reg [31:0] data_234;
  reg [31:0] data_235;
  reg [31:0] data_236;
  reg [31:0] data_237;
  reg [31:0] data_238;
  reg [31:0] data_239;
  reg [31:0] data_240;
  reg [31:0] data_241;
  reg [31:0] data_242;
  reg [31:0] data_243;
  reg [31:0] data_244;
  reg [31:0] data_245;
  reg [31:0] data_246;
  reg [31:0] data_247;
  reg [31:0] data_248;
  reg [31:0] data_249;
  reg [31:0] data_250;
  reg [31:0] data_251;
  reg [31:0] data_252;
  reg [31:0] data_253;
  reg [31:0] data_254;
  reg [31:0] data_255;
  reg [31:0] data_256;
  reg [31:0] data_257;
  reg [31:0] data_258;
  reg [31:0] data_259;
  reg [31:0] data_260;
  reg [31:0] data_261;
  reg [31:0] data_262;
  reg [31:0] data_263;
  reg [31:0] data_264;
  reg [31:0] data_265;
  reg [31:0] data_266;
  reg [31:0] data_267;
  reg [31:0] data_268;
  reg [31:0] data_269;
  reg [31:0] data_270;
  reg [31:0] data_271;
  reg [31:0] data_272;
  reg [31:0] data_273;
  reg [31:0] data_274;
  reg [31:0] data_275;
  reg [31:0] data_276;
  reg [31:0] data_277;
  reg [31:0] data_278;
  reg [31:0] data_279;
  reg [31:0] data_280;
  reg [31:0] data_281;
  reg [31:0] data_282;
  reg [31:0] data_283;
  reg [31:0] data_284;
  reg [31:0] data_285;
  reg [31:0] data_286;
  reg [31:0] data_287;
  reg [31:0] data_288;
  reg [31:0] data_289;
  reg [31:0] data_290;
  reg [31:0] data_291;
  reg [31:0] data_292;
  reg [31:0] data_293;
  reg [31:0] data_294;
  reg [31:0] data_295;
  reg [31:0] data_296;
  reg [31:0] data_297;
  reg [31:0] data_298;
  reg [31:0] data_299;
  reg [31:0] data_300;
  reg [31:0] data_301;
  reg [31:0] data_302;
  reg [31:0] data_303;
  reg [31:0] data_304;
  reg [31:0] data_305;
  reg [31:0] data_306;
  reg [31:0] data_307;
  reg [31:0] data_308;
  reg [31:0] data_309;
  reg [31:0] data_310;
  reg [31:0] data_311;
  reg [31:0] data_312;
  reg [31:0] data_313;
  reg [31:0] data_314;
  reg [31:0] data_315;
  reg [31:0] data_316;
  reg [31:0] data_317;
  reg [31:0] data_318;
  reg [31:0] data_319;
  reg [31:0] data_320;
  reg [31:0] data_321;
  reg [31:0] data_322;
  reg [31:0] data_323;
  reg [31:0] data_324;
  reg [31:0] data_325;
  reg [31:0] data_326;
  reg [31:0] data_327;
  reg [31:0] data_328;
  reg [31:0] data_329;
  reg [31:0] data_330;
  reg [31:0] data_331;
  reg [31:0] data_332;
  reg [31:0] data_333;
  reg [31:0] data_334;
  reg [31:0] data_335;
  reg [31:0] data_336;
  reg [31:0] data_337;
  reg [31:0] data_338;
  reg [31:0] data_339;
  reg [31:0] data_340;
  reg [31:0] data_341;
  reg [31:0] data_342;
  reg [31:0] data_343;
  reg [31:0] data_344;
  reg [31:0] data_345;
  reg [31:0] data_346;
  reg [31:0] data_347;
  reg [31:0] data_348;
  reg [31:0] data_349;
  reg [31:0] data_350;
  reg [31:0] data_351;
  reg [31:0] data_352;
  reg [31:0] data_353;
  reg [31:0] data_354;
  reg [31:0] data_355;
  reg [31:0] data_356;
  reg [31:0] data_357;
  reg [31:0] data_358;
  reg [31:0] data_359;
  reg [31:0] data_360;
  reg [31:0] data_361;
  reg [31:0] data_362;
  reg [31:0] data_363;
  reg [31:0] data_364;
  reg [31:0] data_365;
  reg [31:0] data_366;
  reg [31:0] data_367;
  reg [31:0] data_368;
  reg [31:0] data_369;
  reg [31:0] data_370;
  reg [31:0] data_371;
  reg [31:0] data_372;
  reg [31:0] data_373;
  reg [31:0] data_374;
  reg [31:0] data_375;
  reg [31:0] data_376;
  reg [31:0] data_377;
  reg [31:0] data_378;
  reg [31:0] data_379;
  reg [31:0] data_380;
  reg [31:0] data_381;
  reg [31:0] data_382;
  reg [31:0] data_383;
  reg [31:0] data_384;
  reg [31:0] data_385;
  reg [31:0] data_386;
  reg [31:0] data_387;
  reg [31:0] data_388;
  reg [31:0] data_389;
  reg [31:0] data_390;
  reg [31:0] data_391;
  reg [31:0] data_392;
  reg [31:0] data_393;
  reg [31:0] data_394;
  reg [31:0] data_395;
  reg [31:0] data_396;
  reg [31:0] data_397;
  reg [31:0] data_398;
  reg [31:0] data_399;
  reg [31:0] data_400;
  reg [31:0] data_401;
  reg [31:0] data_402;
  reg [31:0] data_403;
  reg [31:0] data_404;
  reg [31:0] data_405;
  reg [31:0] data_406;
  reg [31:0] data_407;
  reg [31:0] data_408;
  reg [31:0] data_409;
  reg [31:0] data_410;
  reg [31:0] data_411;
  reg [31:0] data_412;
  reg [31:0] data_413;
  reg [31:0] data_414;
  reg [31:0] data_415;
  reg [31:0] data_416;
  reg [31:0] data_417;
  reg [31:0] data_418;
  reg [31:0] data_419;
  reg [31:0] data_420;
  reg [31:0] data_421;
  reg [31:0] data_422;
  reg [31:0] data_423;
  reg [31:0] data_424;
  reg [31:0] data_425;
  reg [31:0] data_426;
  reg [31:0] data_427;
  reg [31:0] data_428;
  reg [31:0] data_429;
  reg [31:0] data_430;
  reg [31:0] data_431;
  reg [31:0] data_432;
  reg [31:0] data_433;
  reg [31:0] data_434;
  reg [31:0] data_435;
  reg [31:0] data_436;
  reg [31:0] data_437;
  reg [31:0] data_438;
  reg [31:0] data_439;
  reg [31:0] data_440;
  reg [31:0] data_441;
  reg [31:0] data_442;
  reg [31:0] data_443;
  reg [31:0] data_444;
  reg [31:0] data_445;
  reg [31:0] data_446;
  reg [31:0] data_447;
  reg [31:0] data_448;
  reg [31:0] data_449;
  reg [31:0] data_450;
  reg [31:0] data_451;
  reg [31:0] data_452;
  reg [31:0] data_453;
  reg [31:0] data_454;
  reg [31:0] data_455;
  reg [31:0] data_456;
  reg [31:0] data_457;
  reg [31:0] data_458;
  reg [31:0] data_459;
  reg [31:0] data_460;
  reg [31:0] data_461;
  reg [31:0] data_462;
  reg [31:0] data_463;
  reg [31:0] data_464;
  reg [31:0] data_465;
  reg [31:0] data_466;
  reg [31:0] data_467;
  reg [31:0] data_468;
  reg [31:0] data_469;
  reg [31:0] data_470;
  reg [31:0] data_471;
  reg [31:0] data_472;
  reg [31:0] data_473;
  reg [31:0] data_474;
  reg [31:0] data_475;
  reg [31:0] data_476;
  reg [31:0] data_477;
  reg [31:0] data_478;
  reg [31:0] data_479;
  reg [31:0] data_480;
  reg [31:0] data_481;
  reg [31:0] data_482;
  reg [31:0] data_483;
  reg [31:0] data_484;
  reg [31:0] data_485;
  reg [31:0] data_486;
  reg [31:0] data_487;
  reg [31:0] data_488;
  reg [31:0] data_489;
  reg [31:0] data_490;
  reg [31:0] data_491;
  reg [31:0] data_492;
  reg [31:0] data_493;
  reg [31:0] data_494;
  reg [31:0] data_495;
  reg [31:0] data_496;
  reg [31:0] data_497;
  reg [31:0] data_498;
  reg [31:0] data_499;
  reg [31:0] data_500;
  reg [31:0] data_501;
  reg [31:0] data_502;
  reg [31:0] data_503;
  reg [31:0] data_504;
  reg [31:0] data_505;
  reg [31:0] data_506;
  reg [31:0] data_507;
  reg [31:0] data_508;
  reg [31:0] data_509;
  reg [31:0] data_510;
  reg [31:0] data_511;
  reg [31:0] data_512;
  reg [31:0] data_513;
  reg [31:0] data_514;
  reg [31:0] data_515;
  reg [31:0] data_516;
  reg [31:0] data_517;
  reg [31:0] data_518;
  reg [31:0] data_519;
  reg [31:0] data_520;
  reg [31:0] data_521;
  reg [31:0] data_522;
  reg [31:0] data_523;
  reg [31:0] data_524;
  reg [31:0] data_525;
  reg [31:0] data_526;
  reg [31:0] data_527;
  reg [31:0] data_528;
  reg [31:0] data_529;
  reg [31:0] data_530;
  reg [31:0] data_531;
  reg [31:0] data_532;
  reg [31:0] data_533;
  reg [31:0] data_534;
  reg [31:0] data_535;
  reg [31:0] data_536;
  reg [31:0] data_537;
  reg [31:0] data_538;
  reg [31:0] data_539;
  reg [31:0] data_540;
  reg [31:0] data_541;
  reg [31:0] data_542;
  reg [31:0] data_543;
  reg [31:0] data_544;
  reg [31:0] data_545;
  reg [31:0] data_546;
  reg [31:0] data_547;
  reg [31:0] data_548;
  reg [31:0] data_549;
  reg [31:0] data_550;
  reg [31:0] data_551;
  reg [31:0] data_552;
  reg [31:0] data_553;
  reg [31:0] data_554;
  reg [31:0] data_555;
  reg [31:0] data_556;
  reg [31:0] data_557;
  reg [31:0] data_558;
  reg [31:0] data_559;
  reg [31:0] data_560;
  reg [31:0] data_561;
  reg [31:0] data_562;
  reg [31:0] data_563;
  reg [31:0] data_564;
  reg [31:0] data_565;
  reg [31:0] data_566;
  reg [31:0] data_567;
  reg [31:0] data_568;
  reg [31:0] data_569;
  reg [31:0] data_570;
  reg [31:0] data_571;
  reg [31:0] data_572;
  reg [31:0] data_573;
  reg [31:0] data_574;
  reg [31:0] data_575;
  reg [31:0] data_576;
  reg [31:0] data_577;
  reg [31:0] data_578;
  reg [31:0] data_579;
  reg [31:0] data_580;
  reg [31:0] data_581;
  reg [31:0] data_582;
  reg [31:0] data_583;
  reg [31:0] data_584;
  reg [31:0] data_585;
  reg [31:0] data_586;
  reg [31:0] data_587;
  reg [31:0] data_588;
  reg [31:0] data_589;
  reg [31:0] data_590;
  reg [31:0] data_591;
  reg [31:0] data_592;
  reg [31:0] data_593;
  reg [31:0] data_594;
  reg [31:0] data_595;
  reg [31:0] data_596;
  reg [31:0] data_597;
  reg [31:0] data_598;
  reg [31:0] data_599;
  reg [31:0] data_600;
  reg [31:0] data_601;
  reg [31:0] data_602;
  reg [31:0] data_603;
  reg [31:0] data_604;
  reg [31:0] data_605;
  reg [31:0] data_606;
  reg [31:0] data_607;
  reg [31:0] data_608;
  reg [31:0] data_609;
  reg [31:0] data_610;
  reg [31:0] data_611;
  reg [31:0] data_612;
  reg [31:0] data_613;
  reg [31:0] data_614;
  reg [31:0] data_615;
  reg [31:0] data_616;
  reg [31:0] data_617;
  reg [31:0] data_618;
  reg [31:0] data_619;
  reg [31:0] data_620;
  reg [31:0] data_621;
  reg [31:0] data_622;
  reg [31:0] data_623;
  reg [31:0] data_624;
  reg [31:0] data_625;
  reg [31:0] data_626;
  reg [31:0] data_627;
  reg [31:0] data_628;
  reg [31:0] data_629;
  reg [31:0] data_630;
  reg [31:0] data_631;
  reg [31:0] data_632;
  reg [31:0] data_633;
  reg [31:0] data_634;
  reg [31:0] data_635;
  reg [31:0] data_636;
  reg [31:0] data_637;
  reg [31:0] data_638;
  reg [31:0] data_639;
  reg [31:0] data_640;
  reg [31:0] data_641;
  reg [31:0] data_642;
  reg [31:0] data_643;
  reg [31:0] data_644;
  reg [31:0] data_645;
  reg [31:0] data_646;
  reg [31:0] data_647;
  reg [31:0] data_648;
  reg [31:0] data_649;
  reg [31:0] data_650;
  reg [31:0] data_651;
  reg [31:0] data_652;
  reg [31:0] data_653;
  reg [31:0] data_654;
  reg [31:0] data_655;
  reg [31:0] data_656;
  reg [31:0] data_657;
  reg [31:0] data_658;
  reg [31:0] data_659;
  reg [31:0] data_660;
  reg [31:0] data_661;
  reg [31:0] data_662;
  reg [31:0] data_663;
  reg [31:0] data_664;
  reg [31:0] data_665;
  reg [31:0] data_666;
  reg [31:0] data_667;
  reg [31:0] data_668;
  reg [31:0] data_669;
  reg [31:0] data_670;
  reg [31:0] data_671;
  reg [31:0] data_672;
  reg [31:0] data_673;
  reg [31:0] data_674;
  reg [31:0] data_675;
  reg [31:0] data_676;
  reg [31:0] data_677;
  reg [31:0] data_678;
  reg [31:0] data_679;
  reg [31:0] data_680;
  reg [31:0] data_681;
  reg [31:0] data_682;
  reg [31:0] data_683;
  reg [31:0] data_684;
  reg [31:0] data_685;
  reg [31:0] data_686;
  reg [31:0] data_687;
  reg [31:0] data_688;
  reg [31:0] data_689;
  reg [31:0] data_690;
  reg [31:0] data_691;
  reg [31:0] data_692;
  reg [31:0] data_693;
  reg [31:0] data_694;
  reg [31:0] data_695;
  reg [31:0] data_696;
  reg [31:0] data_697;
  reg [31:0] data_698;
  reg [31:0] data_699;
  reg [31:0] data_700;
  reg [31:0] data_701;
  reg [31:0] data_702;
  reg [31:0] data_703;
  reg [31:0] data_704;
  reg [31:0] data_705;
  reg [31:0] data_706;
  reg [31:0] data_707;
  reg [31:0] data_708;
  reg [31:0] data_709;
  reg [31:0] data_710;
  reg [31:0] data_711;
  reg [31:0] data_712;
  reg [31:0] data_713;
  reg [31:0] data_714;
  reg [31:0] data_715;
  reg [31:0] data_716;
  reg [31:0] data_717;
  reg [31:0] data_718;
  reg [31:0] data_719;
  reg [31:0] data_720;
  reg [31:0] data_721;
  reg [31:0] data_722;
  reg [31:0] data_723;
  reg [31:0] data_724;
  reg [31:0] data_725;
  reg [31:0] data_726;
  reg [31:0] data_727;
  reg [31:0] data_728;
  reg [31:0] data_729;
  reg [31:0] data_730;
  reg [31:0] data_731;
  reg [31:0] data_732;
  reg [31:0] data_733;
  reg [31:0] data_734;
  reg [31:0] data_735;
  reg [31:0] data_736;
  reg [31:0] data_737;
  reg [31:0] data_738;
  reg [31:0] data_739;
  reg [31:0] data_740;
  reg [31:0] data_741;
  reg [31:0] data_742;
  reg [31:0] data_743;
  reg [31:0] data_744;
  reg [31:0] data_745;
  reg [31:0] data_746;
  reg [31:0] data_747;
  reg [31:0] data_748;
  reg [31:0] data_749;
  reg [31:0] data_750;
  reg [31:0] data_751;
  reg [31:0] data_752;
  reg [31:0] data_753;
  reg [31:0] data_754;
  reg [31:0] data_755;
  reg [31:0] data_756;
  reg [31:0] data_757;
  reg [31:0] data_758;
  reg [31:0] data_759;
  reg [31:0] data_760;
  reg [31:0] data_761;
  reg [31:0] data_762;
  reg [31:0] data_763;
  reg [31:0] data_764;
  reg [31:0] data_765;
  reg [31:0] data_766;
  reg [31:0] data_767;
  reg [31:0] data_768;
  reg [31:0] data_769;
  reg [31:0] data_770;
  reg [31:0] data_771;
  reg [31:0] data_772;
  reg [31:0] data_773;
  reg [31:0] data_774;
  reg [31:0] data_775;
  reg [31:0] data_776;
  reg [31:0] data_777;
  reg [31:0] data_778;
  reg [31:0] data_779;
  reg [31:0] data_780;
  reg [31:0] data_781;
  reg [31:0] data_782;
  reg [31:0] data_783;
  reg [31:0] data_784;
  reg [31:0] data_785;
  reg [31:0] data_786;
  reg [31:0] data_787;
  reg [31:0] data_788;
  reg [31:0] data_789;
  reg [31:0] data_790;
  reg [31:0] data_791;
  reg [31:0] data_792;
  reg [31:0] data_793;
  reg [31:0] data_794;
  reg [31:0] data_795;
  reg [31:0] data_796;
  reg [31:0] data_797;
  reg [31:0] data_798;
  reg [31:0] data_799;
  reg [31:0] data_800;
  reg [31:0] data_801;
  reg [31:0] data_802;
  reg [31:0] data_803;
  reg [31:0] data_804;
  reg [31:0] data_805;
  reg [31:0] data_806;
  reg [31:0] data_807;
  reg [31:0] data_808;
  reg [31:0] data_809;
  reg [31:0] data_810;
  reg [31:0] data_811;
  reg [31:0] data_812;
  reg [31:0] data_813;
  reg [31:0] data_814;
  reg [31:0] data_815;
  reg [31:0] data_816;
  reg [31:0] data_817;
  reg [31:0] data_818;
  reg [31:0] data_819;
  reg [31:0] data_820;
  reg [31:0] data_821;
  reg [31:0] data_822;
  reg [31:0] data_823;
  reg [31:0] data_824;
  reg [31:0] data_825;
  reg [31:0] data_826;
  reg [31:0] data_827;
  reg [31:0] data_828;
  reg [31:0] data_829;
  reg [31:0] data_830;
  reg [31:0] data_831;
  reg [31:0] data_832;
  reg [31:0] data_833;
  reg [31:0] data_834;
  reg [31:0] data_835;
  reg [31:0] data_836;
  reg [31:0] data_837;
  reg [31:0] data_838;
  reg [31:0] data_839;
  reg [31:0] data_840;
  reg [31:0] data_841;
  reg [31:0] data_842;
  reg [31:0] data_843;
  reg [31:0] data_844;
  reg [31:0] data_845;
  reg [31:0] data_846;
  reg [31:0] data_847;
  reg [31:0] data_848;
  reg [31:0] data_849;
  reg [31:0] data_850;
  reg [31:0] data_851;
  reg [31:0] data_852;
  reg [31:0] data_853;
  reg [31:0] data_854;
  reg [31:0] data_855;
  reg [31:0] data_856;
  reg [31:0] data_857;
  reg [31:0] data_858;
  reg [31:0] data_859;
  reg [31:0] data_860;
  reg [31:0] data_861;
  reg [31:0] data_862;
  reg [31:0] data_863;
  reg [31:0] data_864;
  reg [31:0] data_865;
  reg [31:0] data_866;
  reg [31:0] data_867;
  reg [31:0] data_868;
  reg [31:0] data_869;
  reg [31:0] data_870;
  reg [31:0] data_871;
  reg [31:0] data_872;
  reg [31:0] data_873;
  reg [31:0] data_874;
  reg [31:0] data_875;
  reg [31:0] data_876;
  reg [31:0] data_877;
  reg [31:0] data_878;
  reg [31:0] data_879;
  reg [31:0] data_880;
  reg [31:0] data_881;
  reg [31:0] data_882;
  reg [31:0] data_883;
  reg [31:0] data_884;
  reg [31:0] data_885;
  reg [31:0] data_886;
  reg [31:0] data_887;
  reg [31:0] data_888;
  reg [31:0] data_889;
  reg [31:0] data_890;
  reg [31:0] data_891;
  reg [31:0] data_892;
  reg [31:0] data_893;
  reg [31:0] data_894;
  reg [31:0] data_895;
  reg [31:0] data_896;
  reg [31:0] data_897;
  reg [31:0] data_898;
  reg [31:0] data_899;
  reg [31:0] data_900;
  reg [31:0] data_901;
  reg [31:0] data_902;
  reg [31:0] data_903;
  reg [31:0] data_904;
  reg [31:0] data_905;
  reg [31:0] data_906;
  reg [31:0] data_907;
  reg [31:0] data_908;
  reg [31:0] data_909;
  reg [31:0] data_910;
  reg [31:0] data_911;
  reg [31:0] data_912;
  reg [31:0] data_913;
  reg [31:0] data_914;
  reg [31:0] data_915;
  reg [31:0] data_916;
  reg [31:0] data_917;
  reg [31:0] data_918;
  reg [31:0] data_919;
  reg [31:0] data_920;
  reg [31:0] data_921;
  reg [31:0] data_922;
  reg [31:0] data_923;
  reg [31:0] data_924;
  reg [31:0] data_925;
  reg [31:0] data_926;
  reg [31:0] data_927;
  reg [31:0] data_928;
  reg [31:0] data_929;
  reg [31:0] data_930;
  reg [31:0] data_931;
  reg [31:0] data_932;
  reg [31:0] data_933;
  reg [31:0] data_934;
  reg [31:0] data_935;
  reg [31:0] data_936;
  reg [31:0] data_937;
  reg [31:0] data_938;
  reg [31:0] data_939;
  reg [31:0] data_940;
  reg [31:0] data_941;
  reg [31:0] data_942;
  reg [31:0] data_943;
  reg [31:0] data_944;
  reg [31:0] data_945;
  reg [31:0] data_946;
  reg [31:0] data_947;
  reg [31:0] data_948;
  reg [31:0] data_949;
  reg [31:0] data_950;
  reg [31:0] data_951;
  reg [31:0] data_952;
  reg [31:0] data_953;
  reg [31:0] data_954;
  reg [31:0] data_955;
  reg [31:0] data_956;
  reg [31:0] data_957;
  reg [31:0] data_958;
  reg [31:0] data_959;
  reg [31:0] data_960;
  reg [31:0] data_961;
  reg [31:0] data_962;
  reg [31:0] data_963;
  reg [31:0] data_964;
  reg [31:0] data_965;
  reg [31:0] data_966;
  reg [31:0] data_967;
  reg [31:0] data_968;
  reg [31:0] data_969;
  reg [31:0] data_970;
  reg [31:0] data_971;
  reg [31:0] data_972;
  reg [31:0] data_973;
  reg [31:0] data_974;
  reg [31:0] data_975;
  reg [31:0] data_976;
  reg [31:0] data_977;
  reg [31:0] data_978;
  reg [31:0] data_979;
  reg [31:0] data_980;
  reg [31:0] data_981;
  reg [31:0] data_982;
  reg [31:0] data_983;
  reg [31:0] data_984;
  reg [31:0] data_985;
  reg [31:0] data_986;
  reg [31:0] data_987;
  reg [31:0] data_988;
  reg [31:0] data_989;
  reg [31:0] data_990;
  reg [31:0] data_991;
  reg [31:0] data_992;
  reg [31:0] data_993;
  reg [31:0] data_994;
  reg [31:0] data_995;
  reg [31:0] data_996;
  reg [31:0] data_997;
  reg [31:0] data_998;
  reg [31:0] data_999;
  reg [63:0] result;
  wire [63:0] _result_T_1 = $signed(data_0) * $signed(coeffs_0);
  wire [63:0] _result_T_2 = $signed(data_1) * $signed(coeffs_1);
  wire [63:0] _result_T_3 = $signed(data_2) * $signed(coeffs_2);
  wire [63:0] _result_T_4 = $signed(data_3) * $signed(coeffs_3);
  wire [63:0] _result_T_5 = $signed(data_4) * $signed(coeffs_4);
  wire [63:0] _result_T_6 = $signed(data_5) * $signed(coeffs_5);
  wire [63:0] _result_T_7 = $signed(data_6) * $signed(coeffs_6);
  wire [63:0] _result_T_8 = $signed(data_7) * $signed(coeffs_7);
  wire [63:0] _result_T_9 = $signed(data_8) * $signed(coeffs_8);
  wire [63:0] _result_T_10 = $signed(data_9) * $signed(coeffs_9);
  wire [63:0] _result_T_11 = $signed(data_10) * $signed(coeffs_10);
  wire [63:0] _result_T_12 = $signed(data_11) * $signed(coeffs_11);
  wire [63:0] _result_T_13 = $signed(data_12) * $signed(coeffs_12);
  wire [63:0] _result_T_14 = $signed(data_13) * $signed(coeffs_13);
  wire [63:0] _result_T_15 = $signed(data_14) * $signed(coeffs_14);
  wire [63:0] _result_T_16 = $signed(data_15) * $signed(coeffs_15);
  wire [63:0] _result_T_17 = $signed(data_16) * $signed(coeffs_16);
  wire [63:0] _result_T_18 = $signed(data_17) * $signed(coeffs_17);
  wire [63:0] _result_T_19 = $signed(data_18) * $signed(coeffs_18);
  wire [63:0] _result_T_20 = $signed(data_19) * $signed(coeffs_19);
  wire [63:0] _result_T_21 = $signed(data_20) * $signed(coeffs_20);
  wire [63:0] _result_T_22 = $signed(data_21) * $signed(coeffs_21);
  wire [63:0] _result_T_23 = $signed(data_22) * $signed(coeffs_22);
  wire [63:0] _result_T_24 = $signed(data_23) * $signed(coeffs_23);
  wire [63:0] _result_T_25 = $signed(data_24) * $signed(coeffs_24);
  wire [63:0] _result_T_26 = $signed(data_25) * $signed(coeffs_25);
  wire [63:0] _result_T_27 = $signed(data_26) * $signed(coeffs_26);
  wire [63:0] _result_T_28 = $signed(data_27) * $signed(coeffs_27);
  wire [63:0] _result_T_29 = $signed(data_28) * $signed(coeffs_28);
  wire [63:0] _result_T_30 = $signed(data_29) * $signed(coeffs_29);
  wire [63:0] _result_T_31 = $signed(data_30) * $signed(coeffs_30);
  wire [63:0] _result_T_32 = $signed(data_31) * $signed(coeffs_31);
  wire [63:0] _result_T_33 = $signed(data_32) * $signed(coeffs_32);
  wire [63:0] _result_T_34 = $signed(data_33) * $signed(coeffs_33);
  wire [63:0] _result_T_35 = $signed(data_34) * $signed(coeffs_34);
  wire [63:0] _result_T_36 = $signed(data_35) * $signed(coeffs_35);
  wire [63:0] _result_T_37 = $signed(data_36) * $signed(coeffs_36);
  wire [63:0] _result_T_38 = $signed(data_37) * $signed(coeffs_37);
  wire [63:0] _result_T_39 = $signed(data_38) * $signed(coeffs_38);
  wire [63:0] _result_T_40 = $signed(data_39) * $signed(coeffs_39);
  wire [63:0] _result_T_41 = $signed(data_40) * $signed(coeffs_40);
  wire [63:0] _result_T_42 = $signed(data_41) * $signed(coeffs_41);
  wire [63:0] _result_T_43 = $signed(data_42) * $signed(coeffs_42);
  wire [63:0] _result_T_44 = $signed(data_43) * $signed(coeffs_43);
  wire [63:0] _result_T_45 = $signed(data_44) * $signed(coeffs_44);
  wire [63:0] _result_T_46 = $signed(data_45) * $signed(coeffs_45);
  wire [63:0] _result_T_47 = $signed(data_46) * $signed(coeffs_46);
  wire [63:0] _result_T_48 = $signed(data_47) * $signed(coeffs_47);
  wire [63:0] _result_T_49 = $signed(data_48) * $signed(coeffs_48);
  wire [63:0] _result_T_50 = $signed(data_49) * $signed(coeffs_49);
  wire [63:0] _result_T_51 = $signed(data_50) * $signed(coeffs_50);
  wire [63:0] _result_T_52 = $signed(data_51) * $signed(coeffs_51);
  wire [63:0] _result_T_53 = $signed(data_52) * $signed(coeffs_52);
  wire [63:0] _result_T_54 = $signed(data_53) * $signed(coeffs_53);
  wire [63:0] _result_T_55 = $signed(data_54) * $signed(coeffs_54);
  wire [63:0] _result_T_56 = $signed(data_55) * $signed(coeffs_55);
  wire [63:0] _result_T_57 = $signed(data_56) * $signed(coeffs_56);
  wire [63:0] _result_T_58 = $signed(data_57) * $signed(coeffs_57);
  wire [63:0] _result_T_59 = $signed(data_58) * $signed(coeffs_58);
  wire [63:0] _result_T_60 = $signed(data_59) * $signed(coeffs_59);
  wire [63:0] _result_T_61 = $signed(data_60) * $signed(coeffs_60);
  wire [63:0] _result_T_62 = $signed(data_61) * $signed(coeffs_61);
  wire [63:0] _result_T_63 = $signed(data_62) * $signed(coeffs_62);
  wire [63:0] _result_T_64 = $signed(data_63) * $signed(coeffs_63);
  wire [63:0] _result_T_65 = $signed(data_64) * $signed(coeffs_64);
  wire [63:0] _result_T_66 = $signed(data_65) * $signed(coeffs_65);
  wire [63:0] _result_T_67 = $signed(data_66) * $signed(coeffs_66);
  wire [63:0] _result_T_68 = $signed(data_67) * $signed(coeffs_67);
  wire [63:0] _result_T_69 = $signed(data_68) * $signed(coeffs_68);
  wire [63:0] _result_T_70 = $signed(data_69) * $signed(coeffs_69);
  wire [63:0] _result_T_71 = $signed(data_70) * $signed(coeffs_70);
  wire [63:0] _result_T_72 = $signed(data_71) * $signed(coeffs_71);
  wire [63:0] _result_T_73 = $signed(data_72) * $signed(coeffs_72);
  wire [63:0] _result_T_74 = $signed(data_73) * $signed(coeffs_73);
  wire [63:0] _result_T_75 = $signed(data_74) * $signed(coeffs_74);
  wire [63:0] _result_T_76 = $signed(data_75) * $signed(coeffs_75);
  wire [63:0] _result_T_77 = $signed(data_76) * $signed(coeffs_76);
  wire [63:0] _result_T_78 = $signed(data_77) * $signed(coeffs_77);
  wire [63:0] _result_T_79 = $signed(data_78) * $signed(coeffs_78);
  wire [63:0] _result_T_80 = $signed(data_79) * $signed(coeffs_79);
  wire [63:0] _result_T_81 = $signed(data_80) * $signed(coeffs_80);
  wire [63:0] _result_T_82 = $signed(data_81) * $signed(coeffs_81);
  wire [63:0] _result_T_83 = $signed(data_82) * $signed(coeffs_82);
  wire [63:0] _result_T_84 = $signed(data_83) * $signed(coeffs_83);
  wire [63:0] _result_T_85 = $signed(data_84) * $signed(coeffs_84);
  wire [63:0] _result_T_86 = $signed(data_85) * $signed(coeffs_85);
  wire [63:0] _result_T_87 = $signed(data_86) * $signed(coeffs_86);
  wire [63:0] _result_T_88 = $signed(data_87) * $signed(coeffs_87);
  wire [63:0] _result_T_89 = $signed(data_88) * $signed(coeffs_88);
  wire [63:0] _result_T_90 = $signed(data_89) * $signed(coeffs_89);
  wire [63:0] _result_T_91 = $signed(data_90) * $signed(coeffs_90);
  wire [63:0] _result_T_92 = $signed(data_91) * $signed(coeffs_91);
  wire [63:0] _result_T_93 = $signed(data_92) * $signed(coeffs_92);
  wire [63:0] _result_T_94 = $signed(data_93) * $signed(coeffs_93);
  wire [63:0] _result_T_95 = $signed(data_94) * $signed(coeffs_94);
  wire [63:0] _result_T_96 = $signed(data_95) * $signed(coeffs_95);
  wire [63:0] _result_T_97 = $signed(data_96) * $signed(coeffs_96);
  wire [63:0] _result_T_98 = $signed(data_97) * $signed(coeffs_97);
  wire [63:0] _result_T_99 = $signed(data_98) * $signed(coeffs_98);
  wire [63:0] _result_T_100 = $signed(data_99) * $signed(coeffs_99);
  wire [63:0] _result_T_101 = $signed(data_100) * $signed(coeffs_100);
  wire [63:0] _result_T_102 = $signed(data_101) * $signed(coeffs_101);
  wire [63:0] _result_T_103 = $signed(data_102) * $signed(coeffs_102);
  wire [63:0] _result_T_104 = $signed(data_103) * $signed(coeffs_103);
  wire [63:0] _result_T_105 = $signed(data_104) * $signed(coeffs_104);
  wire [63:0] _result_T_106 = $signed(data_105) * $signed(coeffs_105);
  wire [63:0] _result_T_107 = $signed(data_106) * $signed(coeffs_106);
  wire [63:0] _result_T_108 = $signed(data_107) * $signed(coeffs_107);
  wire [63:0] _result_T_109 = $signed(data_108) * $signed(coeffs_108);
  wire [63:0] _result_T_110 = $signed(data_109) * $signed(coeffs_109);
  wire [63:0] _result_T_111 = $signed(data_110) * $signed(coeffs_110);
  wire [63:0] _result_T_112 = $signed(data_111) * $signed(coeffs_111);
  wire [63:0] _result_T_113 = $signed(data_112) * $signed(coeffs_112);
  wire [63:0] _result_T_114 = $signed(data_113) * $signed(coeffs_113);
  wire [63:0] _result_T_115 = $signed(data_114) * $signed(coeffs_114);
  wire [63:0] _result_T_116 = $signed(data_115) * $signed(coeffs_115);
  wire [63:0] _result_T_117 = $signed(data_116) * $signed(coeffs_116);
  wire [63:0] _result_T_118 = $signed(data_117) * $signed(coeffs_117);
  wire [63:0] _result_T_119 = $signed(data_118) * $signed(coeffs_118);
  wire [63:0] _result_T_120 = $signed(data_119) * $signed(coeffs_119);
  wire [63:0] _result_T_121 = $signed(data_120) * $signed(coeffs_120);
  wire [63:0] _result_T_122 = $signed(data_121) * $signed(coeffs_121);
  wire [63:0] _result_T_123 = $signed(data_122) * $signed(coeffs_122);
  wire [63:0] _result_T_124 = $signed(data_123) * $signed(coeffs_123);
  wire [63:0] _result_T_125 = $signed(data_124) * $signed(coeffs_124);
  wire [63:0] _result_T_126 = $signed(data_125) * $signed(coeffs_125);
  wire [63:0] _result_T_127 = $signed(data_126) * $signed(coeffs_126);
  wire [63:0] _result_T_128 = $signed(data_127) * $signed(coeffs_127);
  wire [63:0] _result_T_129 = $signed(data_128) * $signed(coeffs_128);
  wire [63:0] _result_T_130 = $signed(data_129) * $signed(coeffs_129);
  wire [63:0] _result_T_131 = $signed(data_130) * $signed(coeffs_130);
  wire [63:0] _result_T_132 = $signed(data_131) * $signed(coeffs_131);
  wire [63:0] _result_T_133 = $signed(data_132) * $signed(coeffs_132);
  wire [63:0] _result_T_134 = $signed(data_133) * $signed(coeffs_133);
  wire [63:0] _result_T_135 = $signed(data_134) * $signed(coeffs_134);
  wire [63:0] _result_T_136 = $signed(data_135) * $signed(coeffs_135);
  wire [63:0] _result_T_137 = $signed(data_136) * $signed(coeffs_136);
  wire [63:0] _result_T_138 = $signed(data_137) * $signed(coeffs_137);
  wire [63:0] _result_T_139 = $signed(data_138) * $signed(coeffs_138);
  wire [63:0] _result_T_140 = $signed(data_139) * $signed(coeffs_139);
  wire [63:0] _result_T_141 = $signed(data_140) * $signed(coeffs_140);
  wire [63:0] _result_T_142 = $signed(data_141) * $signed(coeffs_141);
  wire [63:0] _result_T_143 = $signed(data_142) * $signed(coeffs_142);
  wire [63:0] _result_T_144 = $signed(data_143) * $signed(coeffs_143);
  wire [63:0] _result_T_145 = $signed(data_144) * $signed(coeffs_144);
  wire [63:0] _result_T_146 = $signed(data_145) * $signed(coeffs_145);
  wire [63:0] _result_T_147 = $signed(data_146) * $signed(coeffs_146);
  wire [63:0] _result_T_148 = $signed(data_147) * $signed(coeffs_147);
  wire [63:0] _result_T_149 = $signed(data_148) * $signed(coeffs_148);
  wire [63:0] _result_T_150 = $signed(data_149) * $signed(coeffs_149);
  wire [63:0] _result_T_151 = $signed(data_150) * $signed(coeffs_150);
  wire [63:0] _result_T_152 = $signed(data_151) * $signed(coeffs_151);
  wire [63:0] _result_T_153 = $signed(data_152) * $signed(coeffs_152);
  wire [63:0] _result_T_154 = $signed(data_153) * $signed(coeffs_153);
  wire [63:0] _result_T_155 = $signed(data_154) * $signed(coeffs_154);
  wire [63:0] _result_T_156 = $signed(data_155) * $signed(coeffs_155);
  wire [63:0] _result_T_157 = $signed(data_156) * $signed(coeffs_156);
  wire [63:0] _result_T_158 = $signed(data_157) * $signed(coeffs_157);
  wire [63:0] _result_T_159 = $signed(data_158) * $signed(coeffs_158);
  wire [63:0] _result_T_160 = $signed(data_159) * $signed(coeffs_159);
  wire [63:0] _result_T_161 = $signed(data_160) * $signed(coeffs_160);
  wire [63:0] _result_T_162 = $signed(data_161) * $signed(coeffs_161);
  wire [63:0] _result_T_163 = $signed(data_162) * $signed(coeffs_162);
  wire [63:0] _result_T_164 = $signed(data_163) * $signed(coeffs_163);
  wire [63:0] _result_T_165 = $signed(data_164) * $signed(coeffs_164);
  wire [63:0] _result_T_166 = $signed(data_165) * $signed(coeffs_165);
  wire [63:0] _result_T_167 = $signed(data_166) * $signed(coeffs_166);
  wire [63:0] _result_T_168 = $signed(data_167) * $signed(coeffs_167);
  wire [63:0] _result_T_169 = $signed(data_168) * $signed(coeffs_168);
  wire [63:0] _result_T_170 = $signed(data_169) * $signed(coeffs_169);
  wire [63:0] _result_T_171 = $signed(data_170) * $signed(coeffs_170);
  wire [63:0] _result_T_172 = $signed(data_171) * $signed(coeffs_171);
  wire [63:0] _result_T_173 = $signed(data_172) * $signed(coeffs_172);
  wire [63:0] _result_T_174 = $signed(data_173) * $signed(coeffs_173);
  wire [63:0] _result_T_175 = $signed(data_174) * $signed(coeffs_174);
  wire [63:0] _result_T_176 = $signed(data_175) * $signed(coeffs_175);
  wire [63:0] _result_T_177 = $signed(data_176) * $signed(coeffs_176);
  wire [63:0] _result_T_178 = $signed(data_177) * $signed(coeffs_177);
  wire [63:0] _result_T_179 = $signed(data_178) * $signed(coeffs_178);
  wire [63:0] _result_T_180 = $signed(data_179) * $signed(coeffs_179);
  wire [63:0] _result_T_181 = $signed(data_180) * $signed(coeffs_180);
  wire [63:0] _result_T_182 = $signed(data_181) * $signed(coeffs_181);
  wire [63:0] _result_T_183 = $signed(data_182) * $signed(coeffs_182);
  wire [63:0] _result_T_184 = $signed(data_183) * $signed(coeffs_183);
  wire [63:0] _result_T_185 = $signed(data_184) * $signed(coeffs_184);
  wire [63:0] _result_T_186 = $signed(data_185) * $signed(coeffs_185);
  wire [63:0] _result_T_187 = $signed(data_186) * $signed(coeffs_186);
  wire [63:0] _result_T_188 = $signed(data_187) * $signed(coeffs_187);
  wire [63:0] _result_T_189 = $signed(data_188) * $signed(coeffs_188);
  wire [63:0] _result_T_190 = $signed(data_189) * $signed(coeffs_189);
  wire [63:0] _result_T_191 = $signed(data_190) * $signed(coeffs_190);
  wire [63:0] _result_T_192 = $signed(data_191) * $signed(coeffs_191);
  wire [63:0] _result_T_193 = $signed(data_192) * $signed(coeffs_192);
  wire [63:0] _result_T_194 = $signed(data_193) * $signed(coeffs_193);
  wire [63:0] _result_T_195 = $signed(data_194) * $signed(coeffs_194);
  wire [63:0] _result_T_196 = $signed(data_195) * $signed(coeffs_195);
  wire [63:0] _result_T_197 = $signed(data_196) * $signed(coeffs_196);
  wire [63:0] _result_T_198 = $signed(data_197) * $signed(coeffs_197);
  wire [63:0] _result_T_199 = $signed(data_198) * $signed(coeffs_198);
  wire [63:0] _result_T_200 = $signed(data_199) * $signed(coeffs_199);
  wire [63:0] _result_T_201 = $signed(data_200) * $signed(coeffs_200);
  wire [63:0] _result_T_202 = $signed(data_201) * $signed(coeffs_201);
  wire [63:0] _result_T_203 = $signed(data_202) * $signed(coeffs_202);
  wire [63:0] _result_T_204 = $signed(data_203) * $signed(coeffs_203);
  wire [63:0] _result_T_205 = $signed(data_204) * $signed(coeffs_204);
  wire [63:0] _result_T_206 = $signed(data_205) * $signed(coeffs_205);
  wire [63:0] _result_T_207 = $signed(data_206) * $signed(coeffs_206);
  wire [63:0] _result_T_208 = $signed(data_207) * $signed(coeffs_207);
  wire [63:0] _result_T_209 = $signed(data_208) * $signed(coeffs_208);
  wire [63:0] _result_T_210 = $signed(data_209) * $signed(coeffs_209);
  wire [63:0] _result_T_211 = $signed(data_210) * $signed(coeffs_210);
  wire [63:0] _result_T_212 = $signed(data_211) * $signed(coeffs_211);
  wire [63:0] _result_T_213 = $signed(data_212) * $signed(coeffs_212);
  wire [63:0] _result_T_214 = $signed(data_213) * $signed(coeffs_213);
  wire [63:0] _result_T_215 = $signed(data_214) * $signed(coeffs_214);
  wire [63:0] _result_T_216 = $signed(data_215) * $signed(coeffs_215);
  wire [63:0] _result_T_217 = $signed(data_216) * $signed(coeffs_216);
  wire [63:0] _result_T_218 = $signed(data_217) * $signed(coeffs_217);
  wire [63:0] _result_T_219 = $signed(data_218) * $signed(coeffs_218);
  wire [63:0] _result_T_220 = $signed(data_219) * $signed(coeffs_219);
  wire [63:0] _result_T_221 = $signed(data_220) * $signed(coeffs_220);
  wire [63:0] _result_T_222 = $signed(data_221) * $signed(coeffs_221);
  wire [63:0] _result_T_223 = $signed(data_222) * $signed(coeffs_222);
  wire [63:0] _result_T_224 = $signed(data_223) * $signed(coeffs_223);
  wire [63:0] _result_T_225 = $signed(data_224) * $signed(coeffs_224);
  wire [63:0] _result_T_226 = $signed(data_225) * $signed(coeffs_225);
  wire [63:0] _result_T_227 = $signed(data_226) * $signed(coeffs_226);
  wire [63:0] _result_T_228 = $signed(data_227) * $signed(coeffs_227);
  wire [63:0] _result_T_229 = $signed(data_228) * $signed(coeffs_228);
  wire [63:0] _result_T_230 = $signed(data_229) * $signed(coeffs_229);
  wire [63:0] _result_T_231 = $signed(data_230) * $signed(coeffs_230);
  wire [63:0] _result_T_232 = $signed(data_231) * $signed(coeffs_231);
  wire [63:0] _result_T_233 = $signed(data_232) * $signed(coeffs_232);
  wire [63:0] _result_T_234 = $signed(data_233) * $signed(coeffs_233);
  wire [63:0] _result_T_235 = $signed(data_234) * $signed(coeffs_234);
  wire [63:0] _result_T_236 = $signed(data_235) * $signed(coeffs_235);
  wire [63:0] _result_T_237 = $signed(data_236) * $signed(coeffs_236);
  wire [63:0] _result_T_238 = $signed(data_237) * $signed(coeffs_237);
  wire [63:0] _result_T_239 = $signed(data_238) * $signed(coeffs_238);
  wire [63:0] _result_T_240 = $signed(data_239) * $signed(coeffs_239);
  wire [63:0] _result_T_241 = $signed(data_240) * $signed(coeffs_240);
  wire [63:0] _result_T_242 = $signed(data_241) * $signed(coeffs_241);
  wire [63:0] _result_T_243 = $signed(data_242) * $signed(coeffs_242);
  wire [63:0] _result_T_244 = $signed(data_243) * $signed(coeffs_243);
  wire [63:0] _result_T_245 = $signed(data_244) * $signed(coeffs_244);
  wire [63:0] _result_T_246 = $signed(data_245) * $signed(coeffs_245);
  wire [63:0] _result_T_247 = $signed(data_246) * $signed(coeffs_246);
  wire [63:0] _result_T_248 = $signed(data_247) * $signed(coeffs_247);
  wire [63:0] _result_T_249 = $signed(data_248) * $signed(coeffs_248);
  wire [63:0] _result_T_250 = $signed(data_249) * $signed(coeffs_249);
  wire [63:0] _result_T_251 = $signed(data_250) * $signed(coeffs_250);
  wire [63:0] _result_T_252 = $signed(data_251) * $signed(coeffs_251);
  wire [63:0] _result_T_253 = $signed(data_252) * $signed(coeffs_252);
  wire [63:0] _result_T_254 = $signed(data_253) * $signed(coeffs_253);
  wire [63:0] _result_T_255 = $signed(data_254) * $signed(coeffs_254);
  wire [63:0] _result_T_256 = $signed(data_255) * $signed(coeffs_255);
  wire [63:0] _result_T_257 = $signed(data_256) * $signed(coeffs_256);
  wire [63:0] _result_T_258 = $signed(data_257) * $signed(coeffs_257);
  wire [63:0] _result_T_259 = $signed(data_258) * $signed(coeffs_258);
  wire [63:0] _result_T_260 = $signed(data_259) * $signed(coeffs_259);
  wire [63:0] _result_T_261 = $signed(data_260) * $signed(coeffs_260);
  wire [63:0] _result_T_262 = $signed(data_261) * $signed(coeffs_261);
  wire [63:0] _result_T_263 = $signed(data_262) * $signed(coeffs_262);
  wire [63:0] _result_T_264 = $signed(data_263) * $signed(coeffs_263);
  wire [63:0] _result_T_265 = $signed(data_264) * $signed(coeffs_264);
  wire [63:0] _result_T_266 = $signed(data_265) * $signed(coeffs_265);
  wire [63:0] _result_T_267 = $signed(data_266) * $signed(coeffs_266);
  wire [63:0] _result_T_268 = $signed(data_267) * $signed(coeffs_267);
  wire [63:0] _result_T_269 = $signed(data_268) * $signed(coeffs_268);
  wire [63:0] _result_T_270 = $signed(data_269) * $signed(coeffs_269);
  wire [63:0] _result_T_271 = $signed(data_270) * $signed(coeffs_270);
  wire [63:0] _result_T_272 = $signed(data_271) * $signed(coeffs_271);
  wire [63:0] _result_T_273 = $signed(data_272) * $signed(coeffs_272);
  wire [63:0] _result_T_274 = $signed(data_273) * $signed(coeffs_273);
  wire [63:0] _result_T_275 = $signed(data_274) * $signed(coeffs_274);
  wire [63:0] _result_T_276 = $signed(data_275) * $signed(coeffs_275);
  wire [63:0] _result_T_277 = $signed(data_276) * $signed(coeffs_276);
  wire [63:0] _result_T_278 = $signed(data_277) * $signed(coeffs_277);
  wire [63:0] _result_T_279 = $signed(data_278) * $signed(coeffs_278);
  wire [63:0] _result_T_280 = $signed(data_279) * $signed(coeffs_279);
  wire [63:0] _result_T_281 = $signed(data_280) * $signed(coeffs_280);
  wire [63:0] _result_T_282 = $signed(data_281) * $signed(coeffs_281);
  wire [63:0] _result_T_283 = $signed(data_282) * $signed(coeffs_282);
  wire [63:0] _result_T_284 = $signed(data_283) * $signed(coeffs_283);
  wire [63:0] _result_T_285 = $signed(data_284) * $signed(coeffs_284);
  wire [63:0] _result_T_286 = $signed(data_285) * $signed(coeffs_285);
  wire [63:0] _result_T_287 = $signed(data_286) * $signed(coeffs_286);
  wire [63:0] _result_T_288 = $signed(data_287) * $signed(coeffs_287);
  wire [63:0] _result_T_289 = $signed(data_288) * $signed(coeffs_288);
  wire [63:0] _result_T_290 = $signed(data_289) * $signed(coeffs_289);
  wire [63:0] _result_T_291 = $signed(data_290) * $signed(coeffs_290);
  wire [63:0] _result_T_292 = $signed(data_291) * $signed(coeffs_291);
  wire [63:0] _result_T_293 = $signed(data_292) * $signed(coeffs_292);
  wire [63:0] _result_T_294 = $signed(data_293) * $signed(coeffs_293);
  wire [63:0] _result_T_295 = $signed(data_294) * $signed(coeffs_294);
  wire [63:0] _result_T_296 = $signed(data_295) * $signed(coeffs_295);
  wire [63:0] _result_T_297 = $signed(data_296) * $signed(coeffs_296);
  wire [63:0] _result_T_298 = $signed(data_297) * $signed(coeffs_297);
  wire [63:0] _result_T_299 = $signed(data_298) * $signed(coeffs_298);
  wire [63:0] _result_T_300 = $signed(data_299) * $signed(coeffs_299);
  wire [63:0] _result_T_301 = $signed(data_300) * $signed(coeffs_300);
  wire [63:0] _result_T_302 = $signed(data_301) * $signed(coeffs_301);
  wire [63:0] _result_T_303 = $signed(data_302) * $signed(coeffs_302);
  wire [63:0] _result_T_304 = $signed(data_303) * $signed(coeffs_303);
  wire [63:0] _result_T_305 = $signed(data_304) * $signed(coeffs_304);
  wire [63:0] _result_T_306 = $signed(data_305) * $signed(coeffs_305);
  wire [63:0] _result_T_307 = $signed(data_306) * $signed(coeffs_306);
  wire [63:0] _result_T_308 = $signed(data_307) * $signed(coeffs_307);
  wire [63:0] _result_T_309 = $signed(data_308) * $signed(coeffs_308);
  wire [63:0] _result_T_310 = $signed(data_309) * $signed(coeffs_309);
  wire [63:0] _result_T_311 = $signed(data_310) * $signed(coeffs_310);
  wire [63:0] _result_T_312 = $signed(data_311) * $signed(coeffs_311);
  wire [63:0] _result_T_313 = $signed(data_312) * $signed(coeffs_312);
  wire [63:0] _result_T_314 = $signed(data_313) * $signed(coeffs_313);
  wire [63:0] _result_T_315 = $signed(data_314) * $signed(coeffs_314);
  wire [63:0] _result_T_316 = $signed(data_315) * $signed(coeffs_315);
  wire [63:0] _result_T_317 = $signed(data_316) * $signed(coeffs_316);
  wire [63:0] _result_T_318 = $signed(data_317) * $signed(coeffs_317);
  wire [63:0] _result_T_319 = $signed(data_318) * $signed(coeffs_318);
  wire [63:0] _result_T_320 = $signed(data_319) * $signed(coeffs_319);
  wire [63:0] _result_T_321 = $signed(data_320) * $signed(coeffs_320);
  wire [63:0] _result_T_322 = $signed(data_321) * $signed(coeffs_321);
  wire [63:0] _result_T_323 = $signed(data_322) * $signed(coeffs_322);
  wire [63:0] _result_T_324 = $signed(data_323) * $signed(coeffs_323);
  wire [63:0] _result_T_325 = $signed(data_324) * $signed(coeffs_324);
  wire [63:0] _result_T_326 = $signed(data_325) * $signed(coeffs_325);
  wire [63:0] _result_T_327 = $signed(data_326) * $signed(coeffs_326);
  wire [63:0] _result_T_328 = $signed(data_327) * $signed(coeffs_327);
  wire [63:0] _result_T_329 = $signed(data_328) * $signed(coeffs_328);
  wire [63:0] _result_T_330 = $signed(data_329) * $signed(coeffs_329);
  wire [63:0] _result_T_331 = $signed(data_330) * $signed(coeffs_330);
  wire [63:0] _result_T_332 = $signed(data_331) * $signed(coeffs_331);
  wire [63:0] _result_T_333 = $signed(data_332) * $signed(coeffs_332);
  wire [63:0] _result_T_334 = $signed(data_333) * $signed(coeffs_333);
  wire [63:0] _result_T_335 = $signed(data_334) * $signed(coeffs_334);
  wire [63:0] _result_T_336 = $signed(data_335) * $signed(coeffs_335);
  wire [63:0] _result_T_337 = $signed(data_336) * $signed(coeffs_336);
  wire [63:0] _result_T_338 = $signed(data_337) * $signed(coeffs_337);
  wire [63:0] _result_T_339 = $signed(data_338) * $signed(coeffs_338);
  wire [63:0] _result_T_340 = $signed(data_339) * $signed(coeffs_339);
  wire [63:0] _result_T_341 = $signed(data_340) * $signed(coeffs_340);
  wire [63:0] _result_T_342 = $signed(data_341) * $signed(coeffs_341);
  wire [63:0] _result_T_343 = $signed(data_342) * $signed(coeffs_342);
  wire [63:0] _result_T_344 = $signed(data_343) * $signed(coeffs_343);
  wire [63:0] _result_T_345 = $signed(data_344) * $signed(coeffs_344);
  wire [63:0] _result_T_346 = $signed(data_345) * $signed(coeffs_345);
  wire [63:0] _result_T_347 = $signed(data_346) * $signed(coeffs_346);
  wire [63:0] _result_T_348 = $signed(data_347) * $signed(coeffs_347);
  wire [63:0] _result_T_349 = $signed(data_348) * $signed(coeffs_348);
  wire [63:0] _result_T_350 = $signed(data_349) * $signed(coeffs_349);
  wire [63:0] _result_T_351 = $signed(data_350) * $signed(coeffs_350);
  wire [63:0] _result_T_352 = $signed(data_351) * $signed(coeffs_351);
  wire [63:0] _result_T_353 = $signed(data_352) * $signed(coeffs_352);
  wire [63:0] _result_T_354 = $signed(data_353) * $signed(coeffs_353);
  wire [63:0] _result_T_355 = $signed(data_354) * $signed(coeffs_354);
  wire [63:0] _result_T_356 = $signed(data_355) * $signed(coeffs_355);
  wire [63:0] _result_T_357 = $signed(data_356) * $signed(coeffs_356);
  wire [63:0] _result_T_358 = $signed(data_357) * $signed(coeffs_357);
  wire [63:0] _result_T_359 = $signed(data_358) * $signed(coeffs_358);
  wire [63:0] _result_T_360 = $signed(data_359) * $signed(coeffs_359);
  wire [63:0] _result_T_361 = $signed(data_360) * $signed(coeffs_360);
  wire [63:0] _result_T_362 = $signed(data_361) * $signed(coeffs_361);
  wire [63:0] _result_T_363 = $signed(data_362) * $signed(coeffs_362);
  wire [63:0] _result_T_364 = $signed(data_363) * $signed(coeffs_363);
  wire [63:0] _result_T_365 = $signed(data_364) * $signed(coeffs_364);
  wire [63:0] _result_T_366 = $signed(data_365) * $signed(coeffs_365);
  wire [63:0] _result_T_367 = $signed(data_366) * $signed(coeffs_366);
  wire [63:0] _result_T_368 = $signed(data_367) * $signed(coeffs_367);
  wire [63:0] _result_T_369 = $signed(data_368) * $signed(coeffs_368);
  wire [63:0] _result_T_370 = $signed(data_369) * $signed(coeffs_369);
  wire [63:0] _result_T_371 = $signed(data_370) * $signed(coeffs_370);
  wire [63:0] _result_T_372 = $signed(data_371) * $signed(coeffs_371);
  wire [63:0] _result_T_373 = $signed(data_372) * $signed(coeffs_372);
  wire [63:0] _result_T_374 = $signed(data_373) * $signed(coeffs_373);
  wire [63:0] _result_T_375 = $signed(data_374) * $signed(coeffs_374);
  wire [63:0] _result_T_376 = $signed(data_375) * $signed(coeffs_375);
  wire [63:0] _result_T_377 = $signed(data_376) * $signed(coeffs_376);
  wire [63:0] _result_T_378 = $signed(data_377) * $signed(coeffs_377);
  wire [63:0] _result_T_379 = $signed(data_378) * $signed(coeffs_378);
  wire [63:0] _result_T_380 = $signed(data_379) * $signed(coeffs_379);
  wire [63:0] _result_T_381 = $signed(data_380) * $signed(coeffs_380);
  wire [63:0] _result_T_382 = $signed(data_381) * $signed(coeffs_381);
  wire [63:0] _result_T_383 = $signed(data_382) * $signed(coeffs_382);
  wire [63:0] _result_T_384 = $signed(data_383) * $signed(coeffs_383);
  wire [63:0] _result_T_385 = $signed(data_384) * $signed(coeffs_384);
  wire [63:0] _result_T_386 = $signed(data_385) * $signed(coeffs_385);
  wire [63:0] _result_T_387 = $signed(data_386) * $signed(coeffs_386);
  wire [63:0] _result_T_388 = $signed(data_387) * $signed(coeffs_387);
  wire [63:0] _result_T_389 = $signed(data_388) * $signed(coeffs_388);
  wire [63:0] _result_T_390 = $signed(data_389) * $signed(coeffs_389);
  wire [63:0] _result_T_391 = $signed(data_390) * $signed(coeffs_390);
  wire [63:0] _result_T_392 = $signed(data_391) * $signed(coeffs_391);
  wire [63:0] _result_T_393 = $signed(data_392) * $signed(coeffs_392);
  wire [63:0] _result_T_394 = $signed(data_393) * $signed(coeffs_393);
  wire [63:0] _result_T_395 = $signed(data_394) * $signed(coeffs_394);
  wire [63:0] _result_T_396 = $signed(data_395) * $signed(coeffs_395);
  wire [63:0] _result_T_397 = $signed(data_396) * $signed(coeffs_396);
  wire [63:0] _result_T_398 = $signed(data_397) * $signed(coeffs_397);
  wire [63:0] _result_T_399 = $signed(data_398) * $signed(coeffs_398);
  wire [63:0] _result_T_400 = $signed(data_399) * $signed(coeffs_399);
  wire [63:0] _result_T_401 = $signed(data_400) * $signed(coeffs_400);
  wire [63:0] _result_T_402 = $signed(data_401) * $signed(coeffs_401);
  wire [63:0] _result_T_403 = $signed(data_402) * $signed(coeffs_402);
  wire [63:0] _result_T_404 = $signed(data_403) * $signed(coeffs_403);
  wire [63:0] _result_T_405 = $signed(data_404) * $signed(coeffs_404);
  wire [63:0] _result_T_406 = $signed(data_405) * $signed(coeffs_405);
  wire [63:0] _result_T_407 = $signed(data_406) * $signed(coeffs_406);
  wire [63:0] _result_T_408 = $signed(data_407) * $signed(coeffs_407);
  wire [63:0] _result_T_409 = $signed(data_408) * $signed(coeffs_408);
  wire [63:0] _result_T_410 = $signed(data_409) * $signed(coeffs_409);
  wire [63:0] _result_T_411 = $signed(data_410) * $signed(coeffs_410);
  wire [63:0] _result_T_412 = $signed(data_411) * $signed(coeffs_411);
  wire [63:0] _result_T_413 = $signed(data_412) * $signed(coeffs_412);
  wire [63:0] _result_T_414 = $signed(data_413) * $signed(coeffs_413);
  wire [63:0] _result_T_415 = $signed(data_414) * $signed(coeffs_414);
  wire [63:0] _result_T_416 = $signed(data_415) * $signed(coeffs_415);
  wire [63:0] _result_T_417 = $signed(data_416) * $signed(coeffs_416);
  wire [63:0] _result_T_418 = $signed(data_417) * $signed(coeffs_417);
  wire [63:0] _result_T_419 = $signed(data_418) * $signed(coeffs_418);
  wire [63:0] _result_T_420 = $signed(data_419) * $signed(coeffs_419);
  wire [63:0] _result_T_421 = $signed(data_420) * $signed(coeffs_420);
  wire [63:0] _result_T_422 = $signed(data_421) * $signed(coeffs_421);
  wire [63:0] _result_T_423 = $signed(data_422) * $signed(coeffs_422);
  wire [63:0] _result_T_424 = $signed(data_423) * $signed(coeffs_423);
  wire [63:0] _result_T_425 = $signed(data_424) * $signed(coeffs_424);
  wire [63:0] _result_T_426 = $signed(data_425) * $signed(coeffs_425);
  wire [63:0] _result_T_427 = $signed(data_426) * $signed(coeffs_426);
  wire [63:0] _result_T_428 = $signed(data_427) * $signed(coeffs_427);
  wire [63:0] _result_T_429 = $signed(data_428) * $signed(coeffs_428);
  wire [63:0] _result_T_430 = $signed(data_429) * $signed(coeffs_429);
  wire [63:0] _result_T_431 = $signed(data_430) * $signed(coeffs_430);
  wire [63:0] _result_T_432 = $signed(data_431) * $signed(coeffs_431);
  wire [63:0] _result_T_433 = $signed(data_432) * $signed(coeffs_432);
  wire [63:0] _result_T_434 = $signed(data_433) * $signed(coeffs_433);
  wire [63:0] _result_T_435 = $signed(data_434) * $signed(coeffs_434);
  wire [63:0] _result_T_436 = $signed(data_435) * $signed(coeffs_435);
  wire [63:0] _result_T_437 = $signed(data_436) * $signed(coeffs_436);
  wire [63:0] _result_T_438 = $signed(data_437) * $signed(coeffs_437);
  wire [63:0] _result_T_439 = $signed(data_438) * $signed(coeffs_438);
  wire [63:0] _result_T_440 = $signed(data_439) * $signed(coeffs_439);
  wire [63:0] _result_T_441 = $signed(data_440) * $signed(coeffs_440);
  wire [63:0] _result_T_442 = $signed(data_441) * $signed(coeffs_441);
  wire [63:0] _result_T_443 = $signed(data_442) * $signed(coeffs_442);
  wire [63:0] _result_T_444 = $signed(data_443) * $signed(coeffs_443);
  wire [63:0] _result_T_445 = $signed(data_444) * $signed(coeffs_444);
  wire [63:0] _result_T_446 = $signed(data_445) * $signed(coeffs_445);
  wire [63:0] _result_T_447 = $signed(data_446) * $signed(coeffs_446);
  wire [63:0] _result_T_448 = $signed(data_447) * $signed(coeffs_447);
  wire [63:0] _result_T_449 = $signed(data_448) * $signed(coeffs_448);
  wire [63:0] _result_T_450 = $signed(data_449) * $signed(coeffs_449);
  wire [63:0] _result_T_451 = $signed(data_450) * $signed(coeffs_450);
  wire [63:0] _result_T_452 = $signed(data_451) * $signed(coeffs_451);
  wire [63:0] _result_T_453 = $signed(data_452) * $signed(coeffs_452);
  wire [63:0] _result_T_454 = $signed(data_453) * $signed(coeffs_453);
  wire [63:0] _result_T_455 = $signed(data_454) * $signed(coeffs_454);
  wire [63:0] _result_T_456 = $signed(data_455) * $signed(coeffs_455);
  wire [63:0] _result_T_457 = $signed(data_456) * $signed(coeffs_456);
  wire [63:0] _result_T_458 = $signed(data_457) * $signed(coeffs_457);
  wire [63:0] _result_T_459 = $signed(data_458) * $signed(coeffs_458);
  wire [63:0] _result_T_460 = $signed(data_459) * $signed(coeffs_459);
  wire [63:0] _result_T_461 = $signed(data_460) * $signed(coeffs_460);
  wire [63:0] _result_T_462 = $signed(data_461) * $signed(coeffs_461);
  wire [63:0] _result_T_463 = $signed(data_462) * $signed(coeffs_462);
  wire [63:0] _result_T_464 = $signed(data_463) * $signed(coeffs_463);
  wire [63:0] _result_T_465 = $signed(data_464) * $signed(coeffs_464);
  wire [63:0] _result_T_466 = $signed(data_465) * $signed(coeffs_465);
  wire [63:0] _result_T_467 = $signed(data_466) * $signed(coeffs_466);
  wire [63:0] _result_T_468 = $signed(data_467) * $signed(coeffs_467);
  wire [63:0] _result_T_469 = $signed(data_468) * $signed(coeffs_468);
  wire [63:0] _result_T_470 = $signed(data_469) * $signed(coeffs_469);
  wire [63:0] _result_T_471 = $signed(data_470) * $signed(coeffs_470);
  wire [63:0] _result_T_472 = $signed(data_471) * $signed(coeffs_471);
  wire [63:0] _result_T_473 = $signed(data_472) * $signed(coeffs_472);
  wire [63:0] _result_T_474 = $signed(data_473) * $signed(coeffs_473);
  wire [63:0] _result_T_475 = $signed(data_474) * $signed(coeffs_474);
  wire [63:0] _result_T_476 = $signed(data_475) * $signed(coeffs_475);
  wire [63:0] _result_T_477 = $signed(data_476) * $signed(coeffs_476);
  wire [63:0] _result_T_478 = $signed(data_477) * $signed(coeffs_477);
  wire [63:0] _result_T_479 = $signed(data_478) * $signed(coeffs_478);
  wire [63:0] _result_T_480 = $signed(data_479) * $signed(coeffs_479);
  wire [63:0] _result_T_481 = $signed(data_480) * $signed(coeffs_480);
  wire [63:0] _result_T_482 = $signed(data_481) * $signed(coeffs_481);
  wire [63:0] _result_T_483 = $signed(data_482) * $signed(coeffs_482);
  wire [63:0] _result_T_484 = $signed(data_483) * $signed(coeffs_483);
  wire [63:0] _result_T_485 = $signed(data_484) * $signed(coeffs_484);
  wire [63:0] _result_T_486 = $signed(data_485) * $signed(coeffs_485);
  wire [63:0] _result_T_487 = $signed(data_486) * $signed(coeffs_486);
  wire [63:0] _result_T_488 = $signed(data_487) * $signed(coeffs_487);
  wire [63:0] _result_T_489 = $signed(data_488) * $signed(coeffs_488);
  wire [63:0] _result_T_490 = $signed(data_489) * $signed(coeffs_489);
  wire [63:0] _result_T_491 = $signed(data_490) * $signed(coeffs_490);
  wire [63:0] _result_T_492 = $signed(data_491) * $signed(coeffs_491);
  wire [63:0] _result_T_493 = $signed(data_492) * $signed(coeffs_492);
  wire [63:0] _result_T_494 = $signed(data_493) * $signed(coeffs_493);
  wire [63:0] _result_T_495 = $signed(data_494) * $signed(coeffs_494);
  wire [63:0] _result_T_496 = $signed(data_495) * $signed(coeffs_495);
  wire [63:0] _result_T_497 = $signed(data_496) * $signed(coeffs_496);
  wire [63:0] _result_T_498 = $signed(data_497) * $signed(coeffs_497);
  wire [63:0] _result_T_499 = $signed(data_498) * $signed(coeffs_498);
  wire [63:0] _result_T_500 = $signed(data_499) * $signed(coeffs_499);
  wire [63:0] _result_T_501 = $signed(data_500) * $signed(coeffs_500);
  wire [63:0] _result_T_502 = $signed(data_501) * $signed(coeffs_501);
  wire [63:0] _result_T_503 = $signed(data_502) * $signed(coeffs_502);
  wire [63:0] _result_T_504 = $signed(data_503) * $signed(coeffs_503);
  wire [63:0] _result_T_505 = $signed(data_504) * $signed(coeffs_504);
  wire [63:0] _result_T_506 = $signed(data_505) * $signed(coeffs_505);
  wire [63:0] _result_T_507 = $signed(data_506) * $signed(coeffs_506);
  wire [63:0] _result_T_508 = $signed(data_507) * $signed(coeffs_507);
  wire [63:0] _result_T_509 = $signed(data_508) * $signed(coeffs_508);
  wire [63:0] _result_T_510 = $signed(data_509) * $signed(coeffs_509);
  wire [63:0] _result_T_511 = $signed(data_510) * $signed(coeffs_510);
  wire [63:0] _result_T_512 = $signed(data_511) * $signed(coeffs_511);
  wire [63:0] _result_T_513 = $signed(data_512) * $signed(coeffs_512);
  wire [63:0] _result_T_514 = $signed(data_513) * $signed(coeffs_513);
  wire [63:0] _result_T_515 = $signed(data_514) * $signed(coeffs_514);
  wire [63:0] _result_T_516 = $signed(data_515) * $signed(coeffs_515);
  wire [63:0] _result_T_517 = $signed(data_516) * $signed(coeffs_516);
  wire [63:0] _result_T_518 = $signed(data_517) * $signed(coeffs_517);
  wire [63:0] _result_T_519 = $signed(data_518) * $signed(coeffs_518);
  wire [63:0] _result_T_520 = $signed(data_519) * $signed(coeffs_519);
  wire [63:0] _result_T_521 = $signed(data_520) * $signed(coeffs_520);
  wire [63:0] _result_T_522 = $signed(data_521) * $signed(coeffs_521);
  wire [63:0] _result_T_523 = $signed(data_522) * $signed(coeffs_522);
  wire [63:0] _result_T_524 = $signed(data_523) * $signed(coeffs_523);
  wire [63:0] _result_T_525 = $signed(data_524) * $signed(coeffs_524);
  wire [63:0] _result_T_526 = $signed(data_525) * $signed(coeffs_525);
  wire [63:0] _result_T_527 = $signed(data_526) * $signed(coeffs_526);
  wire [63:0] _result_T_528 = $signed(data_527) * $signed(coeffs_527);
  wire [63:0] _result_T_529 = $signed(data_528) * $signed(coeffs_528);
  wire [63:0] _result_T_530 = $signed(data_529) * $signed(coeffs_529);
  wire [63:0] _result_T_531 = $signed(data_530) * $signed(coeffs_530);
  wire [63:0] _result_T_532 = $signed(data_531) * $signed(coeffs_531);
  wire [63:0] _result_T_533 = $signed(data_532) * $signed(coeffs_532);
  wire [63:0] _result_T_534 = $signed(data_533) * $signed(coeffs_533);
  wire [63:0] _result_T_535 = $signed(data_534) * $signed(coeffs_534);
  wire [63:0] _result_T_536 = $signed(data_535) * $signed(coeffs_535);
  wire [63:0] _result_T_537 = $signed(data_536) * $signed(coeffs_536);
  wire [63:0] _result_T_538 = $signed(data_537) * $signed(coeffs_537);
  wire [63:0] _result_T_539 = $signed(data_538) * $signed(coeffs_538);
  wire [63:0] _result_T_540 = $signed(data_539) * $signed(coeffs_539);
  wire [63:0] _result_T_541 = $signed(data_540) * $signed(coeffs_540);
  wire [63:0] _result_T_542 = $signed(data_541) * $signed(coeffs_541);
  wire [63:0] _result_T_543 = $signed(data_542) * $signed(coeffs_542);
  wire [63:0] _result_T_544 = $signed(data_543) * $signed(coeffs_543);
  wire [63:0] _result_T_545 = $signed(data_544) * $signed(coeffs_544);
  wire [63:0] _result_T_546 = $signed(data_545) * $signed(coeffs_545);
  wire [63:0] _result_T_547 = $signed(data_546) * $signed(coeffs_546);
  wire [63:0] _result_T_548 = $signed(data_547) * $signed(coeffs_547);
  wire [63:0] _result_T_549 = $signed(data_548) * $signed(coeffs_548);
  wire [63:0] _result_T_550 = $signed(data_549) * $signed(coeffs_549);
  wire [63:0] _result_T_551 = $signed(data_550) * $signed(coeffs_550);
  wire [63:0] _result_T_552 = $signed(data_551) * $signed(coeffs_551);
  wire [63:0] _result_T_553 = $signed(data_552) * $signed(coeffs_552);
  wire [63:0] _result_T_554 = $signed(data_553) * $signed(coeffs_553);
  wire [63:0] _result_T_555 = $signed(data_554) * $signed(coeffs_554);
  wire [63:0] _result_T_556 = $signed(data_555) * $signed(coeffs_555);
  wire [63:0] _result_T_557 = $signed(data_556) * $signed(coeffs_556);
  wire [63:0] _result_T_558 = $signed(data_557) * $signed(coeffs_557);
  wire [63:0] _result_T_559 = $signed(data_558) * $signed(coeffs_558);
  wire [63:0] _result_T_560 = $signed(data_559) * $signed(coeffs_559);
  wire [63:0] _result_T_561 = $signed(data_560) * $signed(coeffs_560);
  wire [63:0] _result_T_562 = $signed(data_561) * $signed(coeffs_561);
  wire [63:0] _result_T_563 = $signed(data_562) * $signed(coeffs_562);
  wire [63:0] _result_T_564 = $signed(data_563) * $signed(coeffs_563);
  wire [63:0] _result_T_565 = $signed(data_564) * $signed(coeffs_564);
  wire [63:0] _result_T_566 = $signed(data_565) * $signed(coeffs_565);
  wire [63:0] _result_T_567 = $signed(data_566) * $signed(coeffs_566);
  wire [63:0] _result_T_568 = $signed(data_567) * $signed(coeffs_567);
  wire [63:0] _result_T_569 = $signed(data_568) * $signed(coeffs_568);
  wire [63:0] _result_T_570 = $signed(data_569) * $signed(coeffs_569);
  wire [63:0] _result_T_571 = $signed(data_570) * $signed(coeffs_570);
  wire [63:0] _result_T_572 = $signed(data_571) * $signed(coeffs_571);
  wire [63:0] _result_T_573 = $signed(data_572) * $signed(coeffs_572);
  wire [63:0] _result_T_574 = $signed(data_573) * $signed(coeffs_573);
  wire [63:0] _result_T_575 = $signed(data_574) * $signed(coeffs_574);
  wire [63:0] _result_T_576 = $signed(data_575) * $signed(coeffs_575);
  wire [63:0] _result_T_577 = $signed(data_576) * $signed(coeffs_576);
  wire [63:0] _result_T_578 = $signed(data_577) * $signed(coeffs_577);
  wire [63:0] _result_T_579 = $signed(data_578) * $signed(coeffs_578);
  wire [63:0] _result_T_580 = $signed(data_579) * $signed(coeffs_579);
  wire [63:0] _result_T_581 = $signed(data_580) * $signed(coeffs_580);
  wire [63:0] _result_T_582 = $signed(data_581) * $signed(coeffs_581);
  wire [63:0] _result_T_583 = $signed(data_582) * $signed(coeffs_582);
  wire [63:0] _result_T_584 = $signed(data_583) * $signed(coeffs_583);
  wire [63:0] _result_T_585 = $signed(data_584) * $signed(coeffs_584);
  wire [63:0] _result_T_586 = $signed(data_585) * $signed(coeffs_585);
  wire [63:0] _result_T_587 = $signed(data_586) * $signed(coeffs_586);
  wire [63:0] _result_T_588 = $signed(data_587) * $signed(coeffs_587);
  wire [63:0] _result_T_589 = $signed(data_588) * $signed(coeffs_588);
  wire [63:0] _result_T_590 = $signed(data_589) * $signed(coeffs_589);
  wire [63:0] _result_T_591 = $signed(data_590) * $signed(coeffs_590);
  wire [63:0] _result_T_592 = $signed(data_591) * $signed(coeffs_591);
  wire [63:0] _result_T_593 = $signed(data_592) * $signed(coeffs_592);
  wire [63:0] _result_T_594 = $signed(data_593) * $signed(coeffs_593);
  wire [63:0] _result_T_595 = $signed(data_594) * $signed(coeffs_594);
  wire [63:0] _result_T_596 = $signed(data_595) * $signed(coeffs_595);
  wire [63:0] _result_T_597 = $signed(data_596) * $signed(coeffs_596);
  wire [63:0] _result_T_598 = $signed(data_597) * $signed(coeffs_597);
  wire [63:0] _result_T_599 = $signed(data_598) * $signed(coeffs_598);
  wire [63:0] _result_T_600 = $signed(data_599) * $signed(coeffs_599);
  wire [63:0] _result_T_601 = $signed(data_600) * $signed(coeffs_600);
  wire [63:0] _result_T_602 = $signed(data_601) * $signed(coeffs_601);
  wire [63:0] _result_T_603 = $signed(data_602) * $signed(coeffs_602);
  wire [63:0] _result_T_604 = $signed(data_603) * $signed(coeffs_603);
  wire [63:0] _result_T_605 = $signed(data_604) * $signed(coeffs_604);
  wire [63:0] _result_T_606 = $signed(data_605) * $signed(coeffs_605);
  wire [63:0] _result_T_607 = $signed(data_606) * $signed(coeffs_606);
  wire [63:0] _result_T_608 = $signed(data_607) * $signed(coeffs_607);
  wire [63:0] _result_T_609 = $signed(data_608) * $signed(coeffs_608);
  wire [63:0] _result_T_610 = $signed(data_609) * $signed(coeffs_609);
  wire [63:0] _result_T_611 = $signed(data_610) * $signed(coeffs_610);
  wire [63:0] _result_T_612 = $signed(data_611) * $signed(coeffs_611);
  wire [63:0] _result_T_613 = $signed(data_612) * $signed(coeffs_612);
  wire [63:0] _result_T_614 = $signed(data_613) * $signed(coeffs_613);
  wire [63:0] _result_T_615 = $signed(data_614) * $signed(coeffs_614);
  wire [63:0] _result_T_616 = $signed(data_615) * $signed(coeffs_615);
  wire [63:0] _result_T_617 = $signed(data_616) * $signed(coeffs_616);
  wire [63:0] _result_T_618 = $signed(data_617) * $signed(coeffs_617);
  wire [63:0] _result_T_619 = $signed(data_618) * $signed(coeffs_618);
  wire [63:0] _result_T_620 = $signed(data_619) * $signed(coeffs_619);
  wire [63:0] _result_T_621 = $signed(data_620) * $signed(coeffs_620);
  wire [63:0] _result_T_622 = $signed(data_621) * $signed(coeffs_621);
  wire [63:0] _result_T_623 = $signed(data_622) * $signed(coeffs_622);
  wire [63:0] _result_T_624 = $signed(data_623) * $signed(coeffs_623);
  wire [63:0] _result_T_625 = $signed(data_624) * $signed(coeffs_624);
  wire [63:0] _result_T_626 = $signed(data_625) * $signed(coeffs_625);
  wire [63:0] _result_T_627 = $signed(data_626) * $signed(coeffs_626);
  wire [63:0] _result_T_628 = $signed(data_627) * $signed(coeffs_627);
  wire [63:0] _result_T_629 = $signed(data_628) * $signed(coeffs_628);
  wire [63:0] _result_T_630 = $signed(data_629) * $signed(coeffs_629);
  wire [63:0] _result_T_631 = $signed(data_630) * $signed(coeffs_630);
  wire [63:0] _result_T_632 = $signed(data_631) * $signed(coeffs_631);
  wire [63:0] _result_T_633 = $signed(data_632) * $signed(coeffs_632);
  wire [63:0] _result_T_634 = $signed(data_633) * $signed(coeffs_633);
  wire [63:0] _result_T_635 = $signed(data_634) * $signed(coeffs_634);
  wire [63:0] _result_T_636 = $signed(data_635) * $signed(coeffs_635);
  wire [63:0] _result_T_637 = $signed(data_636) * $signed(coeffs_636);
  wire [63:0] _result_T_638 = $signed(data_637) * $signed(coeffs_637);
  wire [63:0] _result_T_639 = $signed(data_638) * $signed(coeffs_638);
  wire [63:0] _result_T_640 = $signed(data_639) * $signed(coeffs_639);
  wire [63:0] _result_T_641 = $signed(data_640) * $signed(coeffs_640);
  wire [63:0] _result_T_642 = $signed(data_641) * $signed(coeffs_641);
  wire [63:0] _result_T_643 = $signed(data_642) * $signed(coeffs_642);
  wire [63:0] _result_T_644 = $signed(data_643) * $signed(coeffs_643);
  wire [63:0] _result_T_645 = $signed(data_644) * $signed(coeffs_644);
  wire [63:0] _result_T_646 = $signed(data_645) * $signed(coeffs_645);
  wire [63:0] _result_T_647 = $signed(data_646) * $signed(coeffs_646);
  wire [63:0] _result_T_648 = $signed(data_647) * $signed(coeffs_647);
  wire [63:0] _result_T_649 = $signed(data_648) * $signed(coeffs_648);
  wire [63:0] _result_T_650 = $signed(data_649) * $signed(coeffs_649);
  wire [63:0] _result_T_651 = $signed(data_650) * $signed(coeffs_650);
  wire [63:0] _result_T_652 = $signed(data_651) * $signed(coeffs_651);
  wire [63:0] _result_T_653 = $signed(data_652) * $signed(coeffs_652);
  wire [63:0] _result_T_654 = $signed(data_653) * $signed(coeffs_653);
  wire [63:0] _result_T_655 = $signed(data_654) * $signed(coeffs_654);
  wire [63:0] _result_T_656 = $signed(data_655) * $signed(coeffs_655);
  wire [63:0] _result_T_657 = $signed(data_656) * $signed(coeffs_656);
  wire [63:0] _result_T_658 = $signed(data_657) * $signed(coeffs_657);
  wire [63:0] _result_T_659 = $signed(data_658) * $signed(coeffs_658);
  wire [63:0] _result_T_660 = $signed(data_659) * $signed(coeffs_659);
  wire [63:0] _result_T_661 = $signed(data_660) * $signed(coeffs_660);
  wire [63:0] _result_T_662 = $signed(data_661) * $signed(coeffs_661);
  wire [63:0] _result_T_663 = $signed(data_662) * $signed(coeffs_662);
  wire [63:0] _result_T_664 = $signed(data_663) * $signed(coeffs_663);
  wire [63:0] _result_T_665 = $signed(data_664) * $signed(coeffs_664);
  wire [63:0] _result_T_666 = $signed(data_665) * $signed(coeffs_665);
  wire [63:0] _result_T_667 = $signed(data_666) * $signed(coeffs_666);
  wire [63:0] _result_T_668 = $signed(data_667) * $signed(coeffs_667);
  wire [63:0] _result_T_669 = $signed(data_668) * $signed(coeffs_668);
  wire [63:0] _result_T_670 = $signed(data_669) * $signed(coeffs_669);
  wire [63:0] _result_T_671 = $signed(data_670) * $signed(coeffs_670);
  wire [63:0] _result_T_672 = $signed(data_671) * $signed(coeffs_671);
  wire [63:0] _result_T_673 = $signed(data_672) * $signed(coeffs_672);
  wire [63:0] _result_T_674 = $signed(data_673) * $signed(coeffs_673);
  wire [63:0] _result_T_675 = $signed(data_674) * $signed(coeffs_674);
  wire [63:0] _result_T_676 = $signed(data_675) * $signed(coeffs_675);
  wire [63:0] _result_T_677 = $signed(data_676) * $signed(coeffs_676);
  wire [63:0] _result_T_678 = $signed(data_677) * $signed(coeffs_677);
  wire [63:0] _result_T_679 = $signed(data_678) * $signed(coeffs_678);
  wire [63:0] _result_T_680 = $signed(data_679) * $signed(coeffs_679);
  wire [63:0] _result_T_681 = $signed(data_680) * $signed(coeffs_680);
  wire [63:0] _result_T_682 = $signed(data_681) * $signed(coeffs_681);
  wire [63:0] _result_T_683 = $signed(data_682) * $signed(coeffs_682);
  wire [63:0] _result_T_684 = $signed(data_683) * $signed(coeffs_683);
  wire [63:0] _result_T_685 = $signed(data_684) * $signed(coeffs_684);
  wire [63:0] _result_T_686 = $signed(data_685) * $signed(coeffs_685);
  wire [63:0] _result_T_687 = $signed(data_686) * $signed(coeffs_686);
  wire [63:0] _result_T_688 = $signed(data_687) * $signed(coeffs_687);
  wire [63:0] _result_T_689 = $signed(data_688) * $signed(coeffs_688);
  wire [63:0] _result_T_690 = $signed(data_689) * $signed(coeffs_689);
  wire [63:0] _result_T_691 = $signed(data_690) * $signed(coeffs_690);
  wire [63:0] _result_T_692 = $signed(data_691) * $signed(coeffs_691);
  wire [63:0] _result_T_693 = $signed(data_692) * $signed(coeffs_692);
  wire [63:0] _result_T_694 = $signed(data_693) * $signed(coeffs_693);
  wire [63:0] _result_T_695 = $signed(data_694) * $signed(coeffs_694);
  wire [63:0] _result_T_696 = $signed(data_695) * $signed(coeffs_695);
  wire [63:0] _result_T_697 = $signed(data_696) * $signed(coeffs_696);
  wire [63:0] _result_T_698 = $signed(data_697) * $signed(coeffs_697);
  wire [63:0] _result_T_699 = $signed(data_698) * $signed(coeffs_698);
  wire [63:0] _result_T_700 = $signed(data_699) * $signed(coeffs_699);
  wire [63:0] _result_T_701 = $signed(data_700) * $signed(coeffs_700);
  wire [63:0] _result_T_702 = $signed(data_701) * $signed(coeffs_701);
  wire [63:0] _result_T_703 = $signed(data_702) * $signed(coeffs_702);
  wire [63:0] _result_T_704 = $signed(data_703) * $signed(coeffs_703);
  wire [63:0] _result_T_705 = $signed(data_704) * $signed(coeffs_704);
  wire [63:0] _result_T_706 = $signed(data_705) * $signed(coeffs_705);
  wire [63:0] _result_T_707 = $signed(data_706) * $signed(coeffs_706);
  wire [63:0] _result_T_708 = $signed(data_707) * $signed(coeffs_707);
  wire [63:0] _result_T_709 = $signed(data_708) * $signed(coeffs_708);
  wire [63:0] _result_T_710 = $signed(data_709) * $signed(coeffs_709);
  wire [63:0] _result_T_711 = $signed(data_710) * $signed(coeffs_710);
  wire [63:0] _result_T_712 = $signed(data_711) * $signed(coeffs_711);
  wire [63:0] _result_T_713 = $signed(data_712) * $signed(coeffs_712);
  wire [63:0] _result_T_714 = $signed(data_713) * $signed(coeffs_713);
  wire [63:0] _result_T_715 = $signed(data_714) * $signed(coeffs_714);
  wire [63:0] _result_T_716 = $signed(data_715) * $signed(coeffs_715);
  wire [63:0] _result_T_717 = $signed(data_716) * $signed(coeffs_716);
  wire [63:0] _result_T_718 = $signed(data_717) * $signed(coeffs_717);
  wire [63:0] _result_T_719 = $signed(data_718) * $signed(coeffs_718);
  wire [63:0] _result_T_720 = $signed(data_719) * $signed(coeffs_719);
  wire [63:0] _result_T_721 = $signed(data_720) * $signed(coeffs_720);
  wire [63:0] _result_T_722 = $signed(data_721) * $signed(coeffs_721);
  wire [63:0] _result_T_723 = $signed(data_722) * $signed(coeffs_722);
  wire [63:0] _result_T_724 = $signed(data_723) * $signed(coeffs_723);
  wire [63:0] _result_T_725 = $signed(data_724) * $signed(coeffs_724);
  wire [63:0] _result_T_726 = $signed(data_725) * $signed(coeffs_725);
  wire [63:0] _result_T_727 = $signed(data_726) * $signed(coeffs_726);
  wire [63:0] _result_T_728 = $signed(data_727) * $signed(coeffs_727);
  wire [63:0] _result_T_729 = $signed(data_728) * $signed(coeffs_728);
  wire [63:0] _result_T_730 = $signed(data_729) * $signed(coeffs_729);
  wire [63:0] _result_T_731 = $signed(data_730) * $signed(coeffs_730);
  wire [63:0] _result_T_732 = $signed(data_731) * $signed(coeffs_731);
  wire [63:0] _result_T_733 = $signed(data_732) * $signed(coeffs_732);
  wire [63:0] _result_T_734 = $signed(data_733) * $signed(coeffs_733);
  wire [63:0] _result_T_735 = $signed(data_734) * $signed(coeffs_734);
  wire [63:0] _result_T_736 = $signed(data_735) * $signed(coeffs_735);
  wire [63:0] _result_T_737 = $signed(data_736) * $signed(coeffs_736);
  wire [63:0] _result_T_738 = $signed(data_737) * $signed(coeffs_737);
  wire [63:0] _result_T_739 = $signed(data_738) * $signed(coeffs_738);
  wire [63:0] _result_T_740 = $signed(data_739) * $signed(coeffs_739);
  wire [63:0] _result_T_741 = $signed(data_740) * $signed(coeffs_740);
  wire [63:0] _result_T_742 = $signed(data_741) * $signed(coeffs_741);
  wire [63:0] _result_T_743 = $signed(data_742) * $signed(coeffs_742);
  wire [63:0] _result_T_744 = $signed(data_743) * $signed(coeffs_743);
  wire [63:0] _result_T_745 = $signed(data_744) * $signed(coeffs_744);
  wire [63:0] _result_T_746 = $signed(data_745) * $signed(coeffs_745);
  wire [63:0] _result_T_747 = $signed(data_746) * $signed(coeffs_746);
  wire [63:0] _result_T_748 = $signed(data_747) * $signed(coeffs_747);
  wire [63:0] _result_T_749 = $signed(data_748) * $signed(coeffs_748);
  wire [63:0] _result_T_750 = $signed(data_749) * $signed(coeffs_749);
  wire [63:0] _result_T_751 = $signed(data_750) * $signed(coeffs_750);
  wire [63:0] _result_T_752 = $signed(data_751) * $signed(coeffs_751);
  wire [63:0] _result_T_753 = $signed(data_752) * $signed(coeffs_752);
  wire [63:0] _result_T_754 = $signed(data_753) * $signed(coeffs_753);
  wire [63:0] _result_T_755 = $signed(data_754) * $signed(coeffs_754);
  wire [63:0] _result_T_756 = $signed(data_755) * $signed(coeffs_755);
  wire [63:0] _result_T_757 = $signed(data_756) * $signed(coeffs_756);
  wire [63:0] _result_T_758 = $signed(data_757) * $signed(coeffs_757);
  wire [63:0] _result_T_759 = $signed(data_758) * $signed(coeffs_758);
  wire [63:0] _result_T_760 = $signed(data_759) * $signed(coeffs_759);
  wire [63:0] _result_T_761 = $signed(data_760) * $signed(coeffs_760);
  wire [63:0] _result_T_762 = $signed(data_761) * $signed(coeffs_761);
  wire [63:0] _result_T_763 = $signed(data_762) * $signed(coeffs_762);
  wire [63:0] _result_T_764 = $signed(data_763) * $signed(coeffs_763);
  wire [63:0] _result_T_765 = $signed(data_764) * $signed(coeffs_764);
  wire [63:0] _result_T_766 = $signed(data_765) * $signed(coeffs_765);
  wire [63:0] _result_T_767 = $signed(data_766) * $signed(coeffs_766);
  wire [63:0] _result_T_768 = $signed(data_767) * $signed(coeffs_767);
  wire [63:0] _result_T_769 = $signed(data_768) * $signed(coeffs_768);
  wire [63:0] _result_T_770 = $signed(data_769) * $signed(coeffs_769);
  wire [63:0] _result_T_771 = $signed(data_770) * $signed(coeffs_770);
  wire [63:0] _result_T_772 = $signed(data_771) * $signed(coeffs_771);
  wire [63:0] _result_T_773 = $signed(data_772) * $signed(coeffs_772);
  wire [63:0] _result_T_774 = $signed(data_773) * $signed(coeffs_773);
  wire [63:0] _result_T_775 = $signed(data_774) * $signed(coeffs_774);
  wire [63:0] _result_T_776 = $signed(data_775) * $signed(coeffs_775);
  wire [63:0] _result_T_777 = $signed(data_776) * $signed(coeffs_776);
  wire [63:0] _result_T_778 = $signed(data_777) * $signed(coeffs_777);
  wire [63:0] _result_T_779 = $signed(data_778) * $signed(coeffs_778);
  wire [63:0] _result_T_780 = $signed(data_779) * $signed(coeffs_779);
  wire [63:0] _result_T_781 = $signed(data_780) * $signed(coeffs_780);
  wire [63:0] _result_T_782 = $signed(data_781) * $signed(coeffs_781);
  wire [63:0] _result_T_783 = $signed(data_782) * $signed(coeffs_782);
  wire [63:0] _result_T_784 = $signed(data_783) * $signed(coeffs_783);
  wire [63:0] _result_T_785 = $signed(data_784) * $signed(coeffs_784);
  wire [63:0] _result_T_786 = $signed(data_785) * $signed(coeffs_785);
  wire [63:0] _result_T_787 = $signed(data_786) * $signed(coeffs_786);
  wire [63:0] _result_T_788 = $signed(data_787) * $signed(coeffs_787);
  wire [63:0] _result_T_789 = $signed(data_788) * $signed(coeffs_788);
  wire [63:0] _result_T_790 = $signed(data_789) * $signed(coeffs_789);
  wire [63:0] _result_T_791 = $signed(data_790) * $signed(coeffs_790);
  wire [63:0] _result_T_792 = $signed(data_791) * $signed(coeffs_791);
  wire [63:0] _result_T_793 = $signed(data_792) * $signed(coeffs_792);
  wire [63:0] _result_T_794 = $signed(data_793) * $signed(coeffs_793);
  wire [63:0] _result_T_795 = $signed(data_794) * $signed(coeffs_794);
  wire [63:0] _result_T_796 = $signed(data_795) * $signed(coeffs_795);
  wire [63:0] _result_T_797 = $signed(data_796) * $signed(coeffs_796);
  wire [63:0] _result_T_798 = $signed(data_797) * $signed(coeffs_797);
  wire [63:0] _result_T_799 = $signed(data_798) * $signed(coeffs_798);
  wire [63:0] _result_T_800 = $signed(data_799) * $signed(coeffs_799);
  wire [63:0] _result_T_801 = $signed(data_800) * $signed(coeffs_800);
  wire [63:0] _result_T_802 = $signed(data_801) * $signed(coeffs_801);
  wire [63:0] _result_T_803 = $signed(data_802) * $signed(coeffs_802);
  wire [63:0] _result_T_804 = $signed(data_803) * $signed(coeffs_803);
  wire [63:0] _result_T_805 = $signed(data_804) * $signed(coeffs_804);
  wire [63:0] _result_T_806 = $signed(data_805) * $signed(coeffs_805);
  wire [63:0] _result_T_807 = $signed(data_806) * $signed(coeffs_806);
  wire [63:0] _result_T_808 = $signed(data_807) * $signed(coeffs_807);
  wire [63:0] _result_T_809 = $signed(data_808) * $signed(coeffs_808);
  wire [63:0] _result_T_810 = $signed(data_809) * $signed(coeffs_809);
  wire [63:0] _result_T_811 = $signed(data_810) * $signed(coeffs_810);
  wire [63:0] _result_T_812 = $signed(data_811) * $signed(coeffs_811);
  wire [63:0] _result_T_813 = $signed(data_812) * $signed(coeffs_812);
  wire [63:0] _result_T_814 = $signed(data_813) * $signed(coeffs_813);
  wire [63:0] _result_T_815 = $signed(data_814) * $signed(coeffs_814);
  wire [63:0] _result_T_816 = $signed(data_815) * $signed(coeffs_815);
  wire [63:0] _result_T_817 = $signed(data_816) * $signed(coeffs_816);
  wire [63:0] _result_T_818 = $signed(data_817) * $signed(coeffs_817);
  wire [63:0] _result_T_819 = $signed(data_818) * $signed(coeffs_818);
  wire [63:0] _result_T_820 = $signed(data_819) * $signed(coeffs_819);
  wire [63:0] _result_T_821 = $signed(data_820) * $signed(coeffs_820);
  wire [63:0] _result_T_822 = $signed(data_821) * $signed(coeffs_821);
  wire [63:0] _result_T_823 = $signed(data_822) * $signed(coeffs_822);
  wire [63:0] _result_T_824 = $signed(data_823) * $signed(coeffs_823);
  wire [63:0] _result_T_825 = $signed(data_824) * $signed(coeffs_824);
  wire [63:0] _result_T_826 = $signed(data_825) * $signed(coeffs_825);
  wire [63:0] _result_T_827 = $signed(data_826) * $signed(coeffs_826);
  wire [63:0] _result_T_828 = $signed(data_827) * $signed(coeffs_827);
  wire [63:0] _result_T_829 = $signed(data_828) * $signed(coeffs_828);
  wire [63:0] _result_T_830 = $signed(data_829) * $signed(coeffs_829);
  wire [63:0] _result_T_831 = $signed(data_830) * $signed(coeffs_830);
  wire [63:0] _result_T_832 = $signed(data_831) * $signed(coeffs_831);
  wire [63:0] _result_T_833 = $signed(data_832) * $signed(coeffs_832);
  wire [63:0] _result_T_834 = $signed(data_833) * $signed(coeffs_833);
  wire [63:0] _result_T_835 = $signed(data_834) * $signed(coeffs_834);
  wire [63:0] _result_T_836 = $signed(data_835) * $signed(coeffs_835);
  wire [63:0] _result_T_837 = $signed(data_836) * $signed(coeffs_836);
  wire [63:0] _result_T_838 = $signed(data_837) * $signed(coeffs_837);
  wire [63:0] _result_T_839 = $signed(data_838) * $signed(coeffs_838);
  wire [63:0] _result_T_840 = $signed(data_839) * $signed(coeffs_839);
  wire [63:0] _result_T_841 = $signed(data_840) * $signed(coeffs_840);
  wire [63:0] _result_T_842 = $signed(data_841) * $signed(coeffs_841);
  wire [63:0] _result_T_843 = $signed(data_842) * $signed(coeffs_842);
  wire [63:0] _result_T_844 = $signed(data_843) * $signed(coeffs_843);
  wire [63:0] _result_T_845 = $signed(data_844) * $signed(coeffs_844);
  wire [63:0] _result_T_846 = $signed(data_845) * $signed(coeffs_845);
  wire [63:0] _result_T_847 = $signed(data_846) * $signed(coeffs_846);
  wire [63:0] _result_T_848 = $signed(data_847) * $signed(coeffs_847);
  wire [63:0] _result_T_849 = $signed(data_848) * $signed(coeffs_848);
  wire [63:0] _result_T_850 = $signed(data_849) * $signed(coeffs_849);
  wire [63:0] _result_T_851 = $signed(data_850) * $signed(coeffs_850);
  wire [63:0] _result_T_852 = $signed(data_851) * $signed(coeffs_851);
  wire [63:0] _result_T_853 = $signed(data_852) * $signed(coeffs_852);
  wire [63:0] _result_T_854 = $signed(data_853) * $signed(coeffs_853);
  wire [63:0] _result_T_855 = $signed(data_854) * $signed(coeffs_854);
  wire [63:0] _result_T_856 = $signed(data_855) * $signed(coeffs_855);
  wire [63:0] _result_T_857 = $signed(data_856) * $signed(coeffs_856);
  wire [63:0] _result_T_858 = $signed(data_857) * $signed(coeffs_857);
  wire [63:0] _result_T_859 = $signed(data_858) * $signed(coeffs_858);
  wire [63:0] _result_T_860 = $signed(data_859) * $signed(coeffs_859);
  wire [63:0] _result_T_861 = $signed(data_860) * $signed(coeffs_860);
  wire [63:0] _result_T_862 = $signed(data_861) * $signed(coeffs_861);
  wire [63:0] _result_T_863 = $signed(data_862) * $signed(coeffs_862);
  wire [63:0] _result_T_864 = $signed(data_863) * $signed(coeffs_863);
  wire [63:0] _result_T_865 = $signed(data_864) * $signed(coeffs_864);
  wire [63:0] _result_T_866 = $signed(data_865) * $signed(coeffs_865);
  wire [63:0] _result_T_867 = $signed(data_866) * $signed(coeffs_866);
  wire [63:0] _result_T_868 = $signed(data_867) * $signed(coeffs_867);
  wire [63:0] _result_T_869 = $signed(data_868) * $signed(coeffs_868);
  wire [63:0] _result_T_870 = $signed(data_869) * $signed(coeffs_869);
  wire [63:0] _result_T_871 = $signed(data_870) * $signed(coeffs_870);
  wire [63:0] _result_T_872 = $signed(data_871) * $signed(coeffs_871);
  wire [63:0] _result_T_873 = $signed(data_872) * $signed(coeffs_872);
  wire [63:0] _result_T_874 = $signed(data_873) * $signed(coeffs_873);
  wire [63:0] _result_T_875 = $signed(data_874) * $signed(coeffs_874);
  wire [63:0] _result_T_876 = $signed(data_875) * $signed(coeffs_875);
  wire [63:0] _result_T_877 = $signed(data_876) * $signed(coeffs_876);
  wire [63:0] _result_T_878 = $signed(data_877) * $signed(coeffs_877);
  wire [63:0] _result_T_879 = $signed(data_878) * $signed(coeffs_878);
  wire [63:0] _result_T_880 = $signed(data_879) * $signed(coeffs_879);
  wire [63:0] _result_T_881 = $signed(data_880) * $signed(coeffs_880);
  wire [63:0] _result_T_882 = $signed(data_881) * $signed(coeffs_881);
  wire [63:0] _result_T_883 = $signed(data_882) * $signed(coeffs_882);
  wire [63:0] _result_T_884 = $signed(data_883) * $signed(coeffs_883);
  wire [63:0] _result_T_885 = $signed(data_884) * $signed(coeffs_884);
  wire [63:0] _result_T_886 = $signed(data_885) * $signed(coeffs_885);
  wire [63:0] _result_T_887 = $signed(data_886) * $signed(coeffs_886);
  wire [63:0] _result_T_888 = $signed(data_887) * $signed(coeffs_887);
  wire [63:0] _result_T_889 = $signed(data_888) * $signed(coeffs_888);
  wire [63:0] _result_T_890 = $signed(data_889) * $signed(coeffs_889);
  wire [63:0] _result_T_891 = $signed(data_890) * $signed(coeffs_890);
  wire [63:0] _result_T_892 = $signed(data_891) * $signed(coeffs_891);
  wire [63:0] _result_T_893 = $signed(data_892) * $signed(coeffs_892);
  wire [63:0] _result_T_894 = $signed(data_893) * $signed(coeffs_893);
  wire [63:0] _result_T_895 = $signed(data_894) * $signed(coeffs_894);
  wire [63:0] _result_T_896 = $signed(data_895) * $signed(coeffs_895);
  wire [63:0] _result_T_897 = $signed(data_896) * $signed(coeffs_896);
  wire [63:0] _result_T_898 = $signed(data_897) * $signed(coeffs_897);
  wire [63:0] _result_T_899 = $signed(data_898) * $signed(coeffs_898);
  wire [63:0] _result_T_900 = $signed(data_899) * $signed(coeffs_899);
  wire [63:0] _result_T_901 = $signed(data_900) * $signed(coeffs_900);
  wire [63:0] _result_T_902 = $signed(data_901) * $signed(coeffs_901);
  wire [63:0] _result_T_903 = $signed(data_902) * $signed(coeffs_902);
  wire [63:0] _result_T_904 = $signed(data_903) * $signed(coeffs_903);
  wire [63:0] _result_T_905 = $signed(data_904) * $signed(coeffs_904);
  wire [63:0] _result_T_906 = $signed(data_905) * $signed(coeffs_905);
  wire [63:0] _result_T_907 = $signed(data_906) * $signed(coeffs_906);
  wire [63:0] _result_T_908 = $signed(data_907) * $signed(coeffs_907);
  wire [63:0] _result_T_909 = $signed(data_908) * $signed(coeffs_908);
  wire [63:0] _result_T_910 = $signed(data_909) * $signed(coeffs_909);
  wire [63:0] _result_T_911 = $signed(data_910) * $signed(coeffs_910);
  wire [63:0] _result_T_912 = $signed(data_911) * $signed(coeffs_911);
  wire [63:0] _result_T_913 = $signed(data_912) * $signed(coeffs_912);
  wire [63:0] _result_T_914 = $signed(data_913) * $signed(coeffs_913);
  wire [63:0] _result_T_915 = $signed(data_914) * $signed(coeffs_914);
  wire [63:0] _result_T_916 = $signed(data_915) * $signed(coeffs_915);
  wire [63:0] _result_T_917 = $signed(data_916) * $signed(coeffs_916);
  wire [63:0] _result_T_918 = $signed(data_917) * $signed(coeffs_917);
  wire [63:0] _result_T_919 = $signed(data_918) * $signed(coeffs_918);
  wire [63:0] _result_T_920 = $signed(data_919) * $signed(coeffs_919);
  wire [63:0] _result_T_921 = $signed(data_920) * $signed(coeffs_920);
  wire [63:0] _result_T_922 = $signed(data_921) * $signed(coeffs_921);
  wire [63:0] _result_T_923 = $signed(data_922) * $signed(coeffs_922);
  wire [63:0] _result_T_924 = $signed(data_923) * $signed(coeffs_923);
  wire [63:0] _result_T_925 = $signed(data_924) * $signed(coeffs_924);
  wire [63:0] _result_T_926 = $signed(data_925) * $signed(coeffs_925);
  wire [63:0] _result_T_927 = $signed(data_926) * $signed(coeffs_926);
  wire [63:0] _result_T_928 = $signed(data_927) * $signed(coeffs_927);
  wire [63:0] _result_T_929 = $signed(data_928) * $signed(coeffs_928);
  wire [63:0] _result_T_930 = $signed(data_929) * $signed(coeffs_929);
  wire [63:0] _result_T_931 = $signed(data_930) * $signed(coeffs_930);
  wire [63:0] _result_T_932 = $signed(data_931) * $signed(coeffs_931);
  wire [63:0] _result_T_933 = $signed(data_932) * $signed(coeffs_932);
  wire [63:0] _result_T_934 = $signed(data_933) * $signed(coeffs_933);
  wire [63:0] _result_T_935 = $signed(data_934) * $signed(coeffs_934);
  wire [63:0] _result_T_936 = $signed(data_935) * $signed(coeffs_935);
  wire [63:0] _result_T_937 = $signed(data_936) * $signed(coeffs_936);
  wire [63:0] _result_T_938 = $signed(data_937) * $signed(coeffs_937);
  wire [63:0] _result_T_939 = $signed(data_938) * $signed(coeffs_938);
  wire [63:0] _result_T_940 = $signed(data_939) * $signed(coeffs_939);
  wire [63:0] _result_T_941 = $signed(data_940) * $signed(coeffs_940);
  wire [63:0] _result_T_942 = $signed(data_941) * $signed(coeffs_941);
  wire [63:0] _result_T_943 = $signed(data_942) * $signed(coeffs_942);
  wire [63:0] _result_T_944 = $signed(data_943) * $signed(coeffs_943);
  wire [63:0] _result_T_945 = $signed(data_944) * $signed(coeffs_944);
  wire [63:0] _result_T_946 = $signed(data_945) * $signed(coeffs_945);
  wire [63:0] _result_T_947 = $signed(data_946) * $signed(coeffs_946);
  wire [63:0] _result_T_948 = $signed(data_947) * $signed(coeffs_947);
  wire [63:0] _result_T_949 = $signed(data_948) * $signed(coeffs_948);
  wire [63:0] _result_T_950 = $signed(data_949) * $signed(coeffs_949);
  wire [63:0] _result_T_951 = $signed(data_950) * $signed(coeffs_950);
  wire [63:0] _result_T_952 = $signed(data_951) * $signed(coeffs_951);
  wire [63:0] _result_T_953 = $signed(data_952) * $signed(coeffs_952);
  wire [63:0] _result_T_954 = $signed(data_953) * $signed(coeffs_953);
  wire [63:0] _result_T_955 = $signed(data_954) * $signed(coeffs_954);
  wire [63:0] _result_T_956 = $signed(data_955) * $signed(coeffs_955);
  wire [63:0] _result_T_957 = $signed(data_956) * $signed(coeffs_956);
  wire [63:0] _result_T_958 = $signed(data_957) * $signed(coeffs_957);
  wire [63:0] _result_T_959 = $signed(data_958) * $signed(coeffs_958);
  wire [63:0] _result_T_960 = $signed(data_959) * $signed(coeffs_959);
  wire [63:0] _result_T_961 = $signed(data_960) * $signed(coeffs_960);
  wire [63:0] _result_T_962 = $signed(data_961) * $signed(coeffs_961);
  wire [63:0] _result_T_963 = $signed(data_962) * $signed(coeffs_962);
  wire [63:0] _result_T_964 = $signed(data_963) * $signed(coeffs_963);
  wire [63:0] _result_T_965 = $signed(data_964) * $signed(coeffs_964);
  wire [63:0] _result_T_966 = $signed(data_965) * $signed(coeffs_965);
  wire [63:0] _result_T_967 = $signed(data_966) * $signed(coeffs_966);
  wire [63:0] _result_T_968 = $signed(data_967) * $signed(coeffs_967);
  wire [63:0] _result_T_969 = $signed(data_968) * $signed(coeffs_968);
  wire [63:0] _result_T_970 = $signed(data_969) * $signed(coeffs_969);
  wire [63:0] _result_T_971 = $signed(data_970) * $signed(coeffs_970);
  wire [63:0] _result_T_972 = $signed(data_971) * $signed(coeffs_971);
  wire [63:0] _result_T_973 = $signed(data_972) * $signed(coeffs_972);
  wire [63:0] _result_T_974 = $signed(data_973) * $signed(coeffs_973);
  wire [63:0] _result_T_975 = $signed(data_974) * $signed(coeffs_974);
  wire [63:0] _result_T_976 = $signed(data_975) * $signed(coeffs_975);
  wire [63:0] _result_T_977 = $signed(data_976) * $signed(coeffs_976);
  wire [63:0] _result_T_978 = $signed(data_977) * $signed(coeffs_977);
  wire [63:0] _result_T_979 = $signed(data_978) * $signed(coeffs_978);
  wire [63:0] _result_T_980 = $signed(data_979) * $signed(coeffs_979);
  wire [63:0] _result_T_981 = $signed(data_980) * $signed(coeffs_980);
  wire [63:0] _result_T_982 = $signed(data_981) * $signed(coeffs_981);
  wire [63:0] _result_T_983 = $signed(data_982) * $signed(coeffs_982);
  wire [63:0] _result_T_984 = $signed(data_983) * $signed(coeffs_983);
  wire [63:0] _result_T_985 = $signed(data_984) * $signed(coeffs_984);
  wire [63:0] _result_T_986 = $signed(data_985) * $signed(coeffs_985);
  wire [63:0] _result_T_987 = $signed(data_986) * $signed(coeffs_986);
  wire [63:0] _result_T_988 = $signed(data_987) * $signed(coeffs_987);
  wire [63:0] _result_T_989 = $signed(data_988) * $signed(coeffs_988);
  wire [63:0] _result_T_990 = $signed(data_989) * $signed(coeffs_989);
  wire [63:0] _result_T_991 = $signed(data_990) * $signed(coeffs_990);
  wire [63:0] _result_T_992 = $signed(data_991) * $signed(coeffs_991);
  wire [63:0] _result_T_993 = $signed(data_992) * $signed(coeffs_992);
  wire [63:0] _result_T_994 = $signed(data_993) * $signed(coeffs_993);
  wire [63:0] _result_T_995 = $signed(data_994) * $signed(coeffs_994);
  wire [63:0] _result_T_996 = $signed(data_995) * $signed(coeffs_995);
  wire [63:0] _result_T_997 = $signed(data_996) * $signed(coeffs_996);
  wire [63:0] _result_T_998 = $signed(data_997) * $signed(coeffs_997);
  wire [63:0] _result_T_999 = $signed(data_998) * $signed(coeffs_998);
  wire [63:0] _result_T_1000 = $signed(data_999) * $signed(coeffs_999);
  wire [63:0] _result_T_1003 = $signed(_result_T_1) + $signed(_result_T_2);
  wire [63:0] _result_T_1006 = $signed(_result_T_1003) + $signed(_result_T_3);
  wire [63:0] _result_T_1009 = $signed(_result_T_1006) + $signed(_result_T_4);
  wire [63:0] _result_T_1012 = $signed(_result_T_1009) + $signed(_result_T_5);
  wire [63:0] _result_T_1015 = $signed(_result_T_1012) + $signed(_result_T_6);
  wire [63:0] _result_T_1018 = $signed(_result_T_1015) + $signed(_result_T_7);
  wire [63:0] _result_T_1021 = $signed(_result_T_1018) + $signed(_result_T_8);
  wire [63:0] _result_T_1024 = $signed(_result_T_1021) + $signed(_result_T_9);
  wire [63:0] _result_T_1027 = $signed(_result_T_1024) + $signed(_result_T_10);
  wire [63:0] _result_T_1030 = $signed(_result_T_1027) + $signed(_result_T_11);
  wire [63:0] _result_T_1033 = $signed(_result_T_1030) + $signed(_result_T_12);
  wire [63:0] _result_T_1036 = $signed(_result_T_1033) + $signed(_result_T_13);
  wire [63:0] _result_T_1039 = $signed(_result_T_1036) + $signed(_result_T_14);
  wire [63:0] _result_T_1042 = $signed(_result_T_1039) + $signed(_result_T_15);
  wire [63:0] _result_T_1045 = $signed(_result_T_1042) + $signed(_result_T_16);
  wire [63:0] _result_T_1048 = $signed(_result_T_1045) + $signed(_result_T_17);
  wire [63:0] _result_T_1051 = $signed(_result_T_1048) + $signed(_result_T_18);
  wire [63:0] _result_T_1054 = $signed(_result_T_1051) + $signed(_result_T_19);
  wire [63:0] _result_T_1057 = $signed(_result_T_1054) + $signed(_result_T_20);
  wire [63:0] _result_T_1060 = $signed(_result_T_1057) + $signed(_result_T_21);
  wire [63:0] _result_T_1063 = $signed(_result_T_1060) + $signed(_result_T_22);
  wire [63:0] _result_T_1066 = $signed(_result_T_1063) + $signed(_result_T_23);
  wire [63:0] _result_T_1069 = $signed(_result_T_1066) + $signed(_result_T_24);
  wire [63:0] _result_T_1072 = $signed(_result_T_1069) + $signed(_result_T_25);
  wire [63:0] _result_T_1075 = $signed(_result_T_1072) + $signed(_result_T_26);
  wire [63:0] _result_T_1078 = $signed(_result_T_1075) + $signed(_result_T_27);
  wire [63:0] _result_T_1081 = $signed(_result_T_1078) + $signed(_result_T_28);
  wire [63:0] _result_T_1084 = $signed(_result_T_1081) + $signed(_result_T_29);
  wire [63:0] _result_T_1087 = $signed(_result_T_1084) + $signed(_result_T_30);
  wire [63:0] _result_T_1090 = $signed(_result_T_1087) + $signed(_result_T_31);
  wire [63:0] _result_T_1093 = $signed(_result_T_1090) + $signed(_result_T_32);
  wire [63:0] _result_T_1096 = $signed(_result_T_1093) + $signed(_result_T_33);
  wire [63:0] _result_T_1099 = $signed(_result_T_1096) + $signed(_result_T_34);
  wire [63:0] _result_T_1102 = $signed(_result_T_1099) + $signed(_result_T_35);
  wire [63:0] _result_T_1105 = $signed(_result_T_1102) + $signed(_result_T_36);
  wire [63:0] _result_T_1108 = $signed(_result_T_1105) + $signed(_result_T_37);
  wire [63:0] _result_T_1111 = $signed(_result_T_1108) + $signed(_result_T_38);
  wire [63:0] _result_T_1114 = $signed(_result_T_1111) + $signed(_result_T_39);
  wire [63:0] _result_T_1117 = $signed(_result_T_1114) + $signed(_result_T_40);
  wire [63:0] _result_T_1120 = $signed(_result_T_1117) + $signed(_result_T_41);
  wire [63:0] _result_T_1123 = $signed(_result_T_1120) + $signed(_result_T_42);
  wire [63:0] _result_T_1126 = $signed(_result_T_1123) + $signed(_result_T_43);
  wire [63:0] _result_T_1129 = $signed(_result_T_1126) + $signed(_result_T_44);
  wire [63:0] _result_T_1132 = $signed(_result_T_1129) + $signed(_result_T_45);
  wire [63:0] _result_T_1135 = $signed(_result_T_1132) + $signed(_result_T_46);
  wire [63:0] _result_T_1138 = $signed(_result_T_1135) + $signed(_result_T_47);
  wire [63:0] _result_T_1141 = $signed(_result_T_1138) + $signed(_result_T_48);
  wire [63:0] _result_T_1144 = $signed(_result_T_1141) + $signed(_result_T_49);
  wire [63:0] _result_T_1147 = $signed(_result_T_1144) + $signed(_result_T_50);
  wire [63:0] _result_T_1150 = $signed(_result_T_1147) + $signed(_result_T_51);
  wire [63:0] _result_T_1153 = $signed(_result_T_1150) + $signed(_result_T_52);
  wire [63:0] _result_T_1156 = $signed(_result_T_1153) + $signed(_result_T_53);
  wire [63:0] _result_T_1159 = $signed(_result_T_1156) + $signed(_result_T_54);
  wire [63:0] _result_T_1162 = $signed(_result_T_1159) + $signed(_result_T_55);
  wire [63:0] _result_T_1165 = $signed(_result_T_1162) + $signed(_result_T_56);
  wire [63:0] _result_T_1168 = $signed(_result_T_1165) + $signed(_result_T_57);
  wire [63:0] _result_T_1171 = $signed(_result_T_1168) + $signed(_result_T_58);
  wire [63:0] _result_T_1174 = $signed(_result_T_1171) + $signed(_result_T_59);
  wire [63:0] _result_T_1177 = $signed(_result_T_1174) + $signed(_result_T_60);
  wire [63:0] _result_T_1180 = $signed(_result_T_1177) + $signed(_result_T_61);
  wire [63:0] _result_T_1183 = $signed(_result_T_1180) + $signed(_result_T_62);
  wire [63:0] _result_T_1186 = $signed(_result_T_1183) + $signed(_result_T_63);
  wire [63:0] _result_T_1189 = $signed(_result_T_1186) + $signed(_result_T_64);
  wire [63:0] _result_T_1192 = $signed(_result_T_1189) + $signed(_result_T_65);
  wire [63:0] _result_T_1195 = $signed(_result_T_1192) + $signed(_result_T_66);
  wire [63:0] _result_T_1198 = $signed(_result_T_1195) + $signed(_result_T_67);
  wire [63:0] _result_T_1201 = $signed(_result_T_1198) + $signed(_result_T_68);
  wire [63:0] _result_T_1204 = $signed(_result_T_1201) + $signed(_result_T_69);
  wire [63:0] _result_T_1207 = $signed(_result_T_1204) + $signed(_result_T_70);
  wire [63:0] _result_T_1210 = $signed(_result_T_1207) + $signed(_result_T_71);
  wire [63:0] _result_T_1213 = $signed(_result_T_1210) + $signed(_result_T_72);
  wire [63:0] _result_T_1216 = $signed(_result_T_1213) + $signed(_result_T_73);
  wire [63:0] _result_T_1219 = $signed(_result_T_1216) + $signed(_result_T_74);
  wire [63:0] _result_T_1222 = $signed(_result_T_1219) + $signed(_result_T_75);
  wire [63:0] _result_T_1225 = $signed(_result_T_1222) + $signed(_result_T_76);
  wire [63:0] _result_T_1228 = $signed(_result_T_1225) + $signed(_result_T_77);
  wire [63:0] _result_T_1231 = $signed(_result_T_1228) + $signed(_result_T_78);
  wire [63:0] _result_T_1234 = $signed(_result_T_1231) + $signed(_result_T_79);
  wire [63:0] _result_T_1237 = $signed(_result_T_1234) + $signed(_result_T_80);
  wire [63:0] _result_T_1240 = $signed(_result_T_1237) + $signed(_result_T_81);
  wire [63:0] _result_T_1243 = $signed(_result_T_1240) + $signed(_result_T_82);
  wire [63:0] _result_T_1246 = $signed(_result_T_1243) + $signed(_result_T_83);
  wire [63:0] _result_T_1249 = $signed(_result_T_1246) + $signed(_result_T_84);
  wire [63:0] _result_T_1252 = $signed(_result_T_1249) + $signed(_result_T_85);
  wire [63:0] _result_T_1255 = $signed(_result_T_1252) + $signed(_result_T_86);
  wire [63:0] _result_T_1258 = $signed(_result_T_1255) + $signed(_result_T_87);
  wire [63:0] _result_T_1261 = $signed(_result_T_1258) + $signed(_result_T_88);
  wire [63:0] _result_T_1264 = $signed(_result_T_1261) + $signed(_result_T_89);
  wire [63:0] _result_T_1267 = $signed(_result_T_1264) + $signed(_result_T_90);
  wire [63:0] _result_T_1270 = $signed(_result_T_1267) + $signed(_result_T_91);
  wire [63:0] _result_T_1273 = $signed(_result_T_1270) + $signed(_result_T_92);
  wire [63:0] _result_T_1276 = $signed(_result_T_1273) + $signed(_result_T_93);
  wire [63:0] _result_T_1279 = $signed(_result_T_1276) + $signed(_result_T_94);
  wire [63:0] _result_T_1282 = $signed(_result_T_1279) + $signed(_result_T_95);
  wire [63:0] _result_T_1285 = $signed(_result_T_1282) + $signed(_result_T_96);
  wire [63:0] _result_T_1288 = $signed(_result_T_1285) + $signed(_result_T_97);
  wire [63:0] _result_T_1291 = $signed(_result_T_1288) + $signed(_result_T_98);
  wire [63:0] _result_T_1294 = $signed(_result_T_1291) + $signed(_result_T_99);
  wire [63:0] _result_T_1297 = $signed(_result_T_1294) + $signed(_result_T_100);
  wire [63:0] _result_T_1300 = $signed(_result_T_1297) + $signed(_result_T_101);
  wire [63:0] _result_T_1303 = $signed(_result_T_1300) + $signed(_result_T_102);
  wire [63:0] _result_T_1306 = $signed(_result_T_1303) + $signed(_result_T_103);
  wire [63:0] _result_T_1309 = $signed(_result_T_1306) + $signed(_result_T_104);
  wire [63:0] _result_T_1312 = $signed(_result_T_1309) + $signed(_result_T_105);
  wire [63:0] _result_T_1315 = $signed(_result_T_1312) + $signed(_result_T_106);
  wire [63:0] _result_T_1318 = $signed(_result_T_1315) + $signed(_result_T_107);
  wire [63:0] _result_T_1321 = $signed(_result_T_1318) + $signed(_result_T_108);
  wire [63:0] _result_T_1324 = $signed(_result_T_1321) + $signed(_result_T_109);
  wire [63:0] _result_T_1327 = $signed(_result_T_1324) + $signed(_result_T_110);
  wire [63:0] _result_T_1330 = $signed(_result_T_1327) + $signed(_result_T_111);
  wire [63:0] _result_T_1333 = $signed(_result_T_1330) + $signed(_result_T_112);
  wire [63:0] _result_T_1336 = $signed(_result_T_1333) + $signed(_result_T_113);
  wire [63:0] _result_T_1339 = $signed(_result_T_1336) + $signed(_result_T_114);
  wire [63:0] _result_T_1342 = $signed(_result_T_1339) + $signed(_result_T_115);
  wire [63:0] _result_T_1345 = $signed(_result_T_1342) + $signed(_result_T_116);
  wire [63:0] _result_T_1348 = $signed(_result_T_1345) + $signed(_result_T_117);
  wire [63:0] _result_T_1351 = $signed(_result_T_1348) + $signed(_result_T_118);
  wire [63:0] _result_T_1354 = $signed(_result_T_1351) + $signed(_result_T_119);
  wire [63:0] _result_T_1357 = $signed(_result_T_1354) + $signed(_result_T_120);
  wire [63:0] _result_T_1360 = $signed(_result_T_1357) + $signed(_result_T_121);
  wire [63:0] _result_T_1363 = $signed(_result_T_1360) + $signed(_result_T_122);
  wire [63:0] _result_T_1366 = $signed(_result_T_1363) + $signed(_result_T_123);
  wire [63:0] _result_T_1369 = $signed(_result_T_1366) + $signed(_result_T_124);
  wire [63:0] _result_T_1372 = $signed(_result_T_1369) + $signed(_result_T_125);
  wire [63:0] _result_T_1375 = $signed(_result_T_1372) + $signed(_result_T_126);
  wire [63:0] _result_T_1378 = $signed(_result_T_1375) + $signed(_result_T_127);
  wire [63:0] _result_T_1381 = $signed(_result_T_1378) + $signed(_result_T_128);
  wire [63:0] _result_T_1384 = $signed(_result_T_1381) + $signed(_result_T_129);
  wire [63:0] _result_T_1387 = $signed(_result_T_1384) + $signed(_result_T_130);
  wire [63:0] _result_T_1390 = $signed(_result_T_1387) + $signed(_result_T_131);
  wire [63:0] _result_T_1393 = $signed(_result_T_1390) + $signed(_result_T_132);
  wire [63:0] _result_T_1396 = $signed(_result_T_1393) + $signed(_result_T_133);
  wire [63:0] _result_T_1399 = $signed(_result_T_1396) + $signed(_result_T_134);
  wire [63:0] _result_T_1402 = $signed(_result_T_1399) + $signed(_result_T_135);
  wire [63:0] _result_T_1405 = $signed(_result_T_1402) + $signed(_result_T_136);
  wire [63:0] _result_T_1408 = $signed(_result_T_1405) + $signed(_result_T_137);
  wire [63:0] _result_T_1411 = $signed(_result_T_1408) + $signed(_result_T_138);
  wire [63:0] _result_T_1414 = $signed(_result_T_1411) + $signed(_result_T_139);
  wire [63:0] _result_T_1417 = $signed(_result_T_1414) + $signed(_result_T_140);
  wire [63:0] _result_T_1420 = $signed(_result_T_1417) + $signed(_result_T_141);
  wire [63:0] _result_T_1423 = $signed(_result_T_1420) + $signed(_result_T_142);
  wire [63:0] _result_T_1426 = $signed(_result_T_1423) + $signed(_result_T_143);
  wire [63:0] _result_T_1429 = $signed(_result_T_1426) + $signed(_result_T_144);
  wire [63:0] _result_T_1432 = $signed(_result_T_1429) + $signed(_result_T_145);
  wire [63:0] _result_T_1435 = $signed(_result_T_1432) + $signed(_result_T_146);
  wire [63:0] _result_T_1438 = $signed(_result_T_1435) + $signed(_result_T_147);
  wire [63:0] _result_T_1441 = $signed(_result_T_1438) + $signed(_result_T_148);
  wire [63:0] _result_T_1444 = $signed(_result_T_1441) + $signed(_result_T_149);
  wire [63:0] _result_T_1447 = $signed(_result_T_1444) + $signed(_result_T_150);
  wire [63:0] _result_T_1450 = $signed(_result_T_1447) + $signed(_result_T_151);
  wire [63:0] _result_T_1453 = $signed(_result_T_1450) + $signed(_result_T_152);
  wire [63:0] _result_T_1456 = $signed(_result_T_1453) + $signed(_result_T_153);
  wire [63:0] _result_T_1459 = $signed(_result_T_1456) + $signed(_result_T_154);
  wire [63:0] _result_T_1462 = $signed(_result_T_1459) + $signed(_result_T_155);
  wire [63:0] _result_T_1465 = $signed(_result_T_1462) + $signed(_result_T_156);
  wire [63:0] _result_T_1468 = $signed(_result_T_1465) + $signed(_result_T_157);
  wire [63:0] _result_T_1471 = $signed(_result_T_1468) + $signed(_result_T_158);
  wire [63:0] _result_T_1474 = $signed(_result_T_1471) + $signed(_result_T_159);
  wire [63:0] _result_T_1477 = $signed(_result_T_1474) + $signed(_result_T_160);
  wire [63:0] _result_T_1480 = $signed(_result_T_1477) + $signed(_result_T_161);
  wire [63:0] _result_T_1483 = $signed(_result_T_1480) + $signed(_result_T_162);
  wire [63:0] _result_T_1486 = $signed(_result_T_1483) + $signed(_result_T_163);
  wire [63:0] _result_T_1489 = $signed(_result_T_1486) + $signed(_result_T_164);
  wire [63:0] _result_T_1492 = $signed(_result_T_1489) + $signed(_result_T_165);
  wire [63:0] _result_T_1495 = $signed(_result_T_1492) + $signed(_result_T_166);
  wire [63:0] _result_T_1498 = $signed(_result_T_1495) + $signed(_result_T_167);
  wire [63:0] _result_T_1501 = $signed(_result_T_1498) + $signed(_result_T_168);
  wire [63:0] _result_T_1504 = $signed(_result_T_1501) + $signed(_result_T_169);
  wire [63:0] _result_T_1507 = $signed(_result_T_1504) + $signed(_result_T_170);
  wire [63:0] _result_T_1510 = $signed(_result_T_1507) + $signed(_result_T_171);
  wire [63:0] _result_T_1513 = $signed(_result_T_1510) + $signed(_result_T_172);
  wire [63:0] _result_T_1516 = $signed(_result_T_1513) + $signed(_result_T_173);
  wire [63:0] _result_T_1519 = $signed(_result_T_1516) + $signed(_result_T_174);
  wire [63:0] _result_T_1522 = $signed(_result_T_1519) + $signed(_result_T_175);
  wire [63:0] _result_T_1525 = $signed(_result_T_1522) + $signed(_result_T_176);
  wire [63:0] _result_T_1528 = $signed(_result_T_1525) + $signed(_result_T_177);
  wire [63:0] _result_T_1531 = $signed(_result_T_1528) + $signed(_result_T_178);
  wire [63:0] _result_T_1534 = $signed(_result_T_1531) + $signed(_result_T_179);
  wire [63:0] _result_T_1537 = $signed(_result_T_1534) + $signed(_result_T_180);
  wire [63:0] _result_T_1540 = $signed(_result_T_1537) + $signed(_result_T_181);
  wire [63:0] _result_T_1543 = $signed(_result_T_1540) + $signed(_result_T_182);
  wire [63:0] _result_T_1546 = $signed(_result_T_1543) + $signed(_result_T_183);
  wire [63:0] _result_T_1549 = $signed(_result_T_1546) + $signed(_result_T_184);
  wire [63:0] _result_T_1552 = $signed(_result_T_1549) + $signed(_result_T_185);
  wire [63:0] _result_T_1555 = $signed(_result_T_1552) + $signed(_result_T_186);
  wire [63:0] _result_T_1558 = $signed(_result_T_1555) + $signed(_result_T_187);
  wire [63:0] _result_T_1561 = $signed(_result_T_1558) + $signed(_result_T_188);
  wire [63:0] _result_T_1564 = $signed(_result_T_1561) + $signed(_result_T_189);
  wire [63:0] _result_T_1567 = $signed(_result_T_1564) + $signed(_result_T_190);
  wire [63:0] _result_T_1570 = $signed(_result_T_1567) + $signed(_result_T_191);
  wire [63:0] _result_T_1573 = $signed(_result_T_1570) + $signed(_result_T_192);
  wire [63:0] _result_T_1576 = $signed(_result_T_1573) + $signed(_result_T_193);
  wire [63:0] _result_T_1579 = $signed(_result_T_1576) + $signed(_result_T_194);
  wire [63:0] _result_T_1582 = $signed(_result_T_1579) + $signed(_result_T_195);
  wire [63:0] _result_T_1585 = $signed(_result_T_1582) + $signed(_result_T_196);
  wire [63:0] _result_T_1588 = $signed(_result_T_1585) + $signed(_result_T_197);
  wire [63:0] _result_T_1591 = $signed(_result_T_1588) + $signed(_result_T_198);
  wire [63:0] _result_T_1594 = $signed(_result_T_1591) + $signed(_result_T_199);
  wire [63:0] _result_T_1597 = $signed(_result_T_1594) + $signed(_result_T_200);
  wire [63:0] _result_T_1600 = $signed(_result_T_1597) + $signed(_result_T_201);
  wire [63:0] _result_T_1603 = $signed(_result_T_1600) + $signed(_result_T_202);
  wire [63:0] _result_T_1606 = $signed(_result_T_1603) + $signed(_result_T_203);
  wire [63:0] _result_T_1609 = $signed(_result_T_1606) + $signed(_result_T_204);
  wire [63:0] _result_T_1612 = $signed(_result_T_1609) + $signed(_result_T_205);
  wire [63:0] _result_T_1615 = $signed(_result_T_1612) + $signed(_result_T_206);
  wire [63:0] _result_T_1618 = $signed(_result_T_1615) + $signed(_result_T_207);
  wire [63:0] _result_T_1621 = $signed(_result_T_1618) + $signed(_result_T_208);
  wire [63:0] _result_T_1624 = $signed(_result_T_1621) + $signed(_result_T_209);
  wire [63:0] _result_T_1627 = $signed(_result_T_1624) + $signed(_result_T_210);
  wire [63:0] _result_T_1630 = $signed(_result_T_1627) + $signed(_result_T_211);
  wire [63:0] _result_T_1633 = $signed(_result_T_1630) + $signed(_result_T_212);
  wire [63:0] _result_T_1636 = $signed(_result_T_1633) + $signed(_result_T_213);
  wire [63:0] _result_T_1639 = $signed(_result_T_1636) + $signed(_result_T_214);
  wire [63:0] _result_T_1642 = $signed(_result_T_1639) + $signed(_result_T_215);
  wire [63:0] _result_T_1645 = $signed(_result_T_1642) + $signed(_result_T_216);
  wire [63:0] _result_T_1648 = $signed(_result_T_1645) + $signed(_result_T_217);
  wire [63:0] _result_T_1651 = $signed(_result_T_1648) + $signed(_result_T_218);
  wire [63:0] _result_T_1654 = $signed(_result_T_1651) + $signed(_result_T_219);
  wire [63:0] _result_T_1657 = $signed(_result_T_1654) + $signed(_result_T_220);
  wire [63:0] _result_T_1660 = $signed(_result_T_1657) + $signed(_result_T_221);
  wire [63:0] _result_T_1663 = $signed(_result_T_1660) + $signed(_result_T_222);
  wire [63:0] _result_T_1666 = $signed(_result_T_1663) + $signed(_result_T_223);
  wire [63:0] _result_T_1669 = $signed(_result_T_1666) + $signed(_result_T_224);
  wire [63:0] _result_T_1672 = $signed(_result_T_1669) + $signed(_result_T_225);
  wire [63:0] _result_T_1675 = $signed(_result_T_1672) + $signed(_result_T_226);
  wire [63:0] _result_T_1678 = $signed(_result_T_1675) + $signed(_result_T_227);
  wire [63:0] _result_T_1681 = $signed(_result_T_1678) + $signed(_result_T_228);
  wire [63:0] _result_T_1684 = $signed(_result_T_1681) + $signed(_result_T_229);
  wire [63:0] _result_T_1687 = $signed(_result_T_1684) + $signed(_result_T_230);
  wire [63:0] _result_T_1690 = $signed(_result_T_1687) + $signed(_result_T_231);
  wire [63:0] _result_T_1693 = $signed(_result_T_1690) + $signed(_result_T_232);
  wire [63:0] _result_T_1696 = $signed(_result_T_1693) + $signed(_result_T_233);
  wire [63:0] _result_T_1699 = $signed(_result_T_1696) + $signed(_result_T_234);
  wire [63:0] _result_T_1702 = $signed(_result_T_1699) + $signed(_result_T_235);
  wire [63:0] _result_T_1705 = $signed(_result_T_1702) + $signed(_result_T_236);
  wire [63:0] _result_T_1708 = $signed(_result_T_1705) + $signed(_result_T_237);
  wire [63:0] _result_T_1711 = $signed(_result_T_1708) + $signed(_result_T_238);
  wire [63:0] _result_T_1714 = $signed(_result_T_1711) + $signed(_result_T_239);
  wire [63:0] _result_T_1717 = $signed(_result_T_1714) + $signed(_result_T_240);
  wire [63:0] _result_T_1720 = $signed(_result_T_1717) + $signed(_result_T_241);
  wire [63:0] _result_T_1723 = $signed(_result_T_1720) + $signed(_result_T_242);
  wire [63:0] _result_T_1726 = $signed(_result_T_1723) + $signed(_result_T_243);
  wire [63:0] _result_T_1729 = $signed(_result_T_1726) + $signed(_result_T_244);
  wire [63:0] _result_T_1732 = $signed(_result_T_1729) + $signed(_result_T_245);
  wire [63:0] _result_T_1735 = $signed(_result_T_1732) + $signed(_result_T_246);
  wire [63:0] _result_T_1738 = $signed(_result_T_1735) + $signed(_result_T_247);
  wire [63:0] _result_T_1741 = $signed(_result_T_1738) + $signed(_result_T_248);
  wire [63:0] _result_T_1744 = $signed(_result_T_1741) + $signed(_result_T_249);
  wire [63:0] _result_T_1747 = $signed(_result_T_1744) + $signed(_result_T_250);
  wire [63:0] _result_T_1750 = $signed(_result_T_1747) + $signed(_result_T_251);
  wire [63:0] _result_T_1753 = $signed(_result_T_1750) + $signed(_result_T_252);
  wire [63:0] _result_T_1756 = $signed(_result_T_1753) + $signed(_result_T_253);
  wire [63:0] _result_T_1759 = $signed(_result_T_1756) + $signed(_result_T_254);
  wire [63:0] _result_T_1762 = $signed(_result_T_1759) + $signed(_result_T_255);
  wire [63:0] _result_T_1765 = $signed(_result_T_1762) + $signed(_result_T_256);
  wire [63:0] _result_T_1768 = $signed(_result_T_1765) + $signed(_result_T_257);
  wire [63:0] _result_T_1771 = $signed(_result_T_1768) + $signed(_result_T_258);
  wire [63:0] _result_T_1774 = $signed(_result_T_1771) + $signed(_result_T_259);
  wire [63:0] _result_T_1777 = $signed(_result_T_1774) + $signed(_result_T_260);
  wire [63:0] _result_T_1780 = $signed(_result_T_1777) + $signed(_result_T_261);
  wire [63:0] _result_T_1783 = $signed(_result_T_1780) + $signed(_result_T_262);
  wire [63:0] _result_T_1786 = $signed(_result_T_1783) + $signed(_result_T_263);
  wire [63:0] _result_T_1789 = $signed(_result_T_1786) + $signed(_result_T_264);
  wire [63:0] _result_T_1792 = $signed(_result_T_1789) + $signed(_result_T_265);
  wire [63:0] _result_T_1795 = $signed(_result_T_1792) + $signed(_result_T_266);
  wire [63:0] _result_T_1798 = $signed(_result_T_1795) + $signed(_result_T_267);
  wire [63:0] _result_T_1801 = $signed(_result_T_1798) + $signed(_result_T_268);
  wire [63:0] _result_T_1804 = $signed(_result_T_1801) + $signed(_result_T_269);
  wire [63:0] _result_T_1807 = $signed(_result_T_1804) + $signed(_result_T_270);
  wire [63:0] _result_T_1810 = $signed(_result_T_1807) + $signed(_result_T_271);
  wire [63:0] _result_T_1813 = $signed(_result_T_1810) + $signed(_result_T_272);
  wire [63:0] _result_T_1816 = $signed(_result_T_1813) + $signed(_result_T_273);
  wire [63:0] _result_T_1819 = $signed(_result_T_1816) + $signed(_result_T_274);
  wire [63:0] _result_T_1822 = $signed(_result_T_1819) + $signed(_result_T_275);
  wire [63:0] _result_T_1825 = $signed(_result_T_1822) + $signed(_result_T_276);
  wire [63:0] _result_T_1828 = $signed(_result_T_1825) + $signed(_result_T_277);
  wire [63:0] _result_T_1831 = $signed(_result_T_1828) + $signed(_result_T_278);
  wire [63:0] _result_T_1834 = $signed(_result_T_1831) + $signed(_result_T_279);
  wire [63:0] _result_T_1837 = $signed(_result_T_1834) + $signed(_result_T_280);
  wire [63:0] _result_T_1840 = $signed(_result_T_1837) + $signed(_result_T_281);
  wire [63:0] _result_T_1843 = $signed(_result_T_1840) + $signed(_result_T_282);
  wire [63:0] _result_T_1846 = $signed(_result_T_1843) + $signed(_result_T_283);
  wire [63:0] _result_T_1849 = $signed(_result_T_1846) + $signed(_result_T_284);
  wire [63:0] _result_T_1852 = $signed(_result_T_1849) + $signed(_result_T_285);
  wire [63:0] _result_T_1855 = $signed(_result_T_1852) + $signed(_result_T_286);
  wire [63:0] _result_T_1858 = $signed(_result_T_1855) + $signed(_result_T_287);
  wire [63:0] _result_T_1861 = $signed(_result_T_1858) + $signed(_result_T_288);
  wire [63:0] _result_T_1864 = $signed(_result_T_1861) + $signed(_result_T_289);
  wire [63:0] _result_T_1867 = $signed(_result_T_1864) + $signed(_result_T_290);
  wire [63:0] _result_T_1870 = $signed(_result_T_1867) + $signed(_result_T_291);
  wire [63:0] _result_T_1873 = $signed(_result_T_1870) + $signed(_result_T_292);
  wire [63:0] _result_T_1876 = $signed(_result_T_1873) + $signed(_result_T_293);
  wire [63:0] _result_T_1879 = $signed(_result_T_1876) + $signed(_result_T_294);
  wire [63:0] _result_T_1882 = $signed(_result_T_1879) + $signed(_result_T_295);
  wire [63:0] _result_T_1885 = $signed(_result_T_1882) + $signed(_result_T_296);
  wire [63:0] _result_T_1888 = $signed(_result_T_1885) + $signed(_result_T_297);
  wire [63:0] _result_T_1891 = $signed(_result_T_1888) + $signed(_result_T_298);
  wire [63:0] _result_T_1894 = $signed(_result_T_1891) + $signed(_result_T_299);
  wire [63:0] _result_T_1897 = $signed(_result_T_1894) + $signed(_result_T_300);
  wire [63:0] _result_T_1900 = $signed(_result_T_1897) + $signed(_result_T_301);
  wire [63:0] _result_T_1903 = $signed(_result_T_1900) + $signed(_result_T_302);
  wire [63:0] _result_T_1906 = $signed(_result_T_1903) + $signed(_result_T_303);
  wire [63:0] _result_T_1909 = $signed(_result_T_1906) + $signed(_result_T_304);
  wire [63:0] _result_T_1912 = $signed(_result_T_1909) + $signed(_result_T_305);
  wire [63:0] _result_T_1915 = $signed(_result_T_1912) + $signed(_result_T_306);
  wire [63:0] _result_T_1918 = $signed(_result_T_1915) + $signed(_result_T_307);
  wire [63:0] _result_T_1921 = $signed(_result_T_1918) + $signed(_result_T_308);
  wire [63:0] _result_T_1924 = $signed(_result_T_1921) + $signed(_result_T_309);
  wire [63:0] _result_T_1927 = $signed(_result_T_1924) + $signed(_result_T_310);
  wire [63:0] _result_T_1930 = $signed(_result_T_1927) + $signed(_result_T_311);
  wire [63:0] _result_T_1933 = $signed(_result_T_1930) + $signed(_result_T_312);
  wire [63:0] _result_T_1936 = $signed(_result_T_1933) + $signed(_result_T_313);
  wire [63:0] _result_T_1939 = $signed(_result_T_1936) + $signed(_result_T_314);
  wire [63:0] _result_T_1942 = $signed(_result_T_1939) + $signed(_result_T_315);
  wire [63:0] _result_T_1945 = $signed(_result_T_1942) + $signed(_result_T_316);
  wire [63:0] _result_T_1948 = $signed(_result_T_1945) + $signed(_result_T_317);
  wire [63:0] _result_T_1951 = $signed(_result_T_1948) + $signed(_result_T_318);
  wire [63:0] _result_T_1954 = $signed(_result_T_1951) + $signed(_result_T_319);
  wire [63:0] _result_T_1957 = $signed(_result_T_1954) + $signed(_result_T_320);
  wire [63:0] _result_T_1960 = $signed(_result_T_1957) + $signed(_result_T_321);
  wire [63:0] _result_T_1963 = $signed(_result_T_1960) + $signed(_result_T_322);
  wire [63:0] _result_T_1966 = $signed(_result_T_1963) + $signed(_result_T_323);
  wire [63:0] _result_T_1969 = $signed(_result_T_1966) + $signed(_result_T_324);
  wire [63:0] _result_T_1972 = $signed(_result_T_1969) + $signed(_result_T_325);
  wire [63:0] _result_T_1975 = $signed(_result_T_1972) + $signed(_result_T_326);
  wire [63:0] _result_T_1978 = $signed(_result_T_1975) + $signed(_result_T_327);
  wire [63:0] _result_T_1981 = $signed(_result_T_1978) + $signed(_result_T_328);
  wire [63:0] _result_T_1984 = $signed(_result_T_1981) + $signed(_result_T_329);
  wire [63:0] _result_T_1987 = $signed(_result_T_1984) + $signed(_result_T_330);
  wire [63:0] _result_T_1990 = $signed(_result_T_1987) + $signed(_result_T_331);
  wire [63:0] _result_T_1993 = $signed(_result_T_1990) + $signed(_result_T_332);
  wire [63:0] _result_T_1996 = $signed(_result_T_1993) + $signed(_result_T_333);
  wire [63:0] _result_T_1999 = $signed(_result_T_1996) + $signed(_result_T_334);
  wire [63:0] _result_T_2002 = $signed(_result_T_1999) + $signed(_result_T_335);
  wire [63:0] _result_T_2005 = $signed(_result_T_2002) + $signed(_result_T_336);
  wire [63:0] _result_T_2008 = $signed(_result_T_2005) + $signed(_result_T_337);
  wire [63:0] _result_T_2011 = $signed(_result_T_2008) + $signed(_result_T_338);
  wire [63:0] _result_T_2014 = $signed(_result_T_2011) + $signed(_result_T_339);
  wire [63:0] _result_T_2017 = $signed(_result_T_2014) + $signed(_result_T_340);
  wire [63:0] _result_T_2020 = $signed(_result_T_2017) + $signed(_result_T_341);
  wire [63:0] _result_T_2023 = $signed(_result_T_2020) + $signed(_result_T_342);
  wire [63:0] _result_T_2026 = $signed(_result_T_2023) + $signed(_result_T_343);
  wire [63:0] _result_T_2029 = $signed(_result_T_2026) + $signed(_result_T_344);
  wire [63:0] _result_T_2032 = $signed(_result_T_2029) + $signed(_result_T_345);
  wire [63:0] _result_T_2035 = $signed(_result_T_2032) + $signed(_result_T_346);
  wire [63:0] _result_T_2038 = $signed(_result_T_2035) + $signed(_result_T_347);
  wire [63:0] _result_T_2041 = $signed(_result_T_2038) + $signed(_result_T_348);
  wire [63:0] _result_T_2044 = $signed(_result_T_2041) + $signed(_result_T_349);
  wire [63:0] _result_T_2047 = $signed(_result_T_2044) + $signed(_result_T_350);
  wire [63:0] _result_T_2050 = $signed(_result_T_2047) + $signed(_result_T_351);
  wire [63:0] _result_T_2053 = $signed(_result_T_2050) + $signed(_result_T_352);
  wire [63:0] _result_T_2056 = $signed(_result_T_2053) + $signed(_result_T_353);
  wire [63:0] _result_T_2059 = $signed(_result_T_2056) + $signed(_result_T_354);
  wire [63:0] _result_T_2062 = $signed(_result_T_2059) + $signed(_result_T_355);
  wire [63:0] _result_T_2065 = $signed(_result_T_2062) + $signed(_result_T_356);
  wire [63:0] _result_T_2068 = $signed(_result_T_2065) + $signed(_result_T_357);
  wire [63:0] _result_T_2071 = $signed(_result_T_2068) + $signed(_result_T_358);
  wire [63:0] _result_T_2074 = $signed(_result_T_2071) + $signed(_result_T_359);
  wire [63:0] _result_T_2077 = $signed(_result_T_2074) + $signed(_result_T_360);
  wire [63:0] _result_T_2080 = $signed(_result_T_2077) + $signed(_result_T_361);
  wire [63:0] _result_T_2083 = $signed(_result_T_2080) + $signed(_result_T_362);
  wire [63:0] _result_T_2086 = $signed(_result_T_2083) + $signed(_result_T_363);
  wire [63:0] _result_T_2089 = $signed(_result_T_2086) + $signed(_result_T_364);
  wire [63:0] _result_T_2092 = $signed(_result_T_2089) + $signed(_result_T_365);
  wire [63:0] _result_T_2095 = $signed(_result_T_2092) + $signed(_result_T_366);
  wire [63:0] _result_T_2098 = $signed(_result_T_2095) + $signed(_result_T_367);
  wire [63:0] _result_T_2101 = $signed(_result_T_2098) + $signed(_result_T_368);
  wire [63:0] _result_T_2104 = $signed(_result_T_2101) + $signed(_result_T_369);
  wire [63:0] _result_T_2107 = $signed(_result_T_2104) + $signed(_result_T_370);
  wire [63:0] _result_T_2110 = $signed(_result_T_2107) + $signed(_result_T_371);
  wire [63:0] _result_T_2113 = $signed(_result_T_2110) + $signed(_result_T_372);
  wire [63:0] _result_T_2116 = $signed(_result_T_2113) + $signed(_result_T_373);
  wire [63:0] _result_T_2119 = $signed(_result_T_2116) + $signed(_result_T_374);
  wire [63:0] _result_T_2122 = $signed(_result_T_2119) + $signed(_result_T_375);
  wire [63:0] _result_T_2125 = $signed(_result_T_2122) + $signed(_result_T_376);
  wire [63:0] _result_T_2128 = $signed(_result_T_2125) + $signed(_result_T_377);
  wire [63:0] _result_T_2131 = $signed(_result_T_2128) + $signed(_result_T_378);
  wire [63:0] _result_T_2134 = $signed(_result_T_2131) + $signed(_result_T_379);
  wire [63:0] _result_T_2137 = $signed(_result_T_2134) + $signed(_result_T_380);
  wire [63:0] _result_T_2140 = $signed(_result_T_2137) + $signed(_result_T_381);
  wire [63:0] _result_T_2143 = $signed(_result_T_2140) + $signed(_result_T_382);
  wire [63:0] _result_T_2146 = $signed(_result_T_2143) + $signed(_result_T_383);
  wire [63:0] _result_T_2149 = $signed(_result_T_2146) + $signed(_result_T_384);
  wire [63:0] _result_T_2152 = $signed(_result_T_2149) + $signed(_result_T_385);
  wire [63:0] _result_T_2155 = $signed(_result_T_2152) + $signed(_result_T_386);
  wire [63:0] _result_T_2158 = $signed(_result_T_2155) + $signed(_result_T_387);
  wire [63:0] _result_T_2161 = $signed(_result_T_2158) + $signed(_result_T_388);
  wire [63:0] _result_T_2164 = $signed(_result_T_2161) + $signed(_result_T_389);
  wire [63:0] _result_T_2167 = $signed(_result_T_2164) + $signed(_result_T_390);
  wire [63:0] _result_T_2170 = $signed(_result_T_2167) + $signed(_result_T_391);
  wire [63:0] _result_T_2173 = $signed(_result_T_2170) + $signed(_result_T_392);
  wire [63:0] _result_T_2176 = $signed(_result_T_2173) + $signed(_result_T_393);
  wire [63:0] _result_T_2179 = $signed(_result_T_2176) + $signed(_result_T_394);
  wire [63:0] _result_T_2182 = $signed(_result_T_2179) + $signed(_result_T_395);
  wire [63:0] _result_T_2185 = $signed(_result_T_2182) + $signed(_result_T_396);
  wire [63:0] _result_T_2188 = $signed(_result_T_2185) + $signed(_result_T_397);
  wire [63:0] _result_T_2191 = $signed(_result_T_2188) + $signed(_result_T_398);
  wire [63:0] _result_T_2194 = $signed(_result_T_2191) + $signed(_result_T_399);
  wire [63:0] _result_T_2197 = $signed(_result_T_2194) + $signed(_result_T_400);
  wire [63:0] _result_T_2200 = $signed(_result_T_2197) + $signed(_result_T_401);
  wire [63:0] _result_T_2203 = $signed(_result_T_2200) + $signed(_result_T_402);
  wire [63:0] _result_T_2206 = $signed(_result_T_2203) + $signed(_result_T_403);
  wire [63:0] _result_T_2209 = $signed(_result_T_2206) + $signed(_result_T_404);
  wire [63:0] _result_T_2212 = $signed(_result_T_2209) + $signed(_result_T_405);
  wire [63:0] _result_T_2215 = $signed(_result_T_2212) + $signed(_result_T_406);
  wire [63:0] _result_T_2218 = $signed(_result_T_2215) + $signed(_result_T_407);
  wire [63:0] _result_T_2221 = $signed(_result_T_2218) + $signed(_result_T_408);
  wire [63:0] _result_T_2224 = $signed(_result_T_2221) + $signed(_result_T_409);
  wire [63:0] _result_T_2227 = $signed(_result_T_2224) + $signed(_result_T_410);
  wire [63:0] _result_T_2230 = $signed(_result_T_2227) + $signed(_result_T_411);
  wire [63:0] _result_T_2233 = $signed(_result_T_2230) + $signed(_result_T_412);
  wire [63:0] _result_T_2236 = $signed(_result_T_2233) + $signed(_result_T_413);
  wire [63:0] _result_T_2239 = $signed(_result_T_2236) + $signed(_result_T_414);
  wire [63:0] _result_T_2242 = $signed(_result_T_2239) + $signed(_result_T_415);
  wire [63:0] _result_T_2245 = $signed(_result_T_2242) + $signed(_result_T_416);
  wire [63:0] _result_T_2248 = $signed(_result_T_2245) + $signed(_result_T_417);
  wire [63:0] _result_T_2251 = $signed(_result_T_2248) + $signed(_result_T_418);
  wire [63:0] _result_T_2254 = $signed(_result_T_2251) + $signed(_result_T_419);
  wire [63:0] _result_T_2257 = $signed(_result_T_2254) + $signed(_result_T_420);
  wire [63:0] _result_T_2260 = $signed(_result_T_2257) + $signed(_result_T_421);
  wire [63:0] _result_T_2263 = $signed(_result_T_2260) + $signed(_result_T_422);
  wire [63:0] _result_T_2266 = $signed(_result_T_2263) + $signed(_result_T_423);
  wire [63:0] _result_T_2269 = $signed(_result_T_2266) + $signed(_result_T_424);
  wire [63:0] _result_T_2272 = $signed(_result_T_2269) + $signed(_result_T_425);
  wire [63:0] _result_T_2275 = $signed(_result_T_2272) + $signed(_result_T_426);
  wire [63:0] _result_T_2278 = $signed(_result_T_2275) + $signed(_result_T_427);
  wire [63:0] _result_T_2281 = $signed(_result_T_2278) + $signed(_result_T_428);
  wire [63:0] _result_T_2284 = $signed(_result_T_2281) + $signed(_result_T_429);
  wire [63:0] _result_T_2287 = $signed(_result_T_2284) + $signed(_result_T_430);
  wire [63:0] _result_T_2290 = $signed(_result_T_2287) + $signed(_result_T_431);
  wire [63:0] _result_T_2293 = $signed(_result_T_2290) + $signed(_result_T_432);
  wire [63:0] _result_T_2296 = $signed(_result_T_2293) + $signed(_result_T_433);
  wire [63:0] _result_T_2299 = $signed(_result_T_2296) + $signed(_result_T_434);
  wire [63:0] _result_T_2302 = $signed(_result_T_2299) + $signed(_result_T_435);
  wire [63:0] _result_T_2305 = $signed(_result_T_2302) + $signed(_result_T_436);
  wire [63:0] _result_T_2308 = $signed(_result_T_2305) + $signed(_result_T_437);
  wire [63:0] _result_T_2311 = $signed(_result_T_2308) + $signed(_result_T_438);
  wire [63:0] _result_T_2314 = $signed(_result_T_2311) + $signed(_result_T_439);
  wire [63:0] _result_T_2317 = $signed(_result_T_2314) + $signed(_result_T_440);
  wire [63:0] _result_T_2320 = $signed(_result_T_2317) + $signed(_result_T_441);
  wire [63:0] _result_T_2323 = $signed(_result_T_2320) + $signed(_result_T_442);
  wire [63:0] _result_T_2326 = $signed(_result_T_2323) + $signed(_result_T_443);
  wire [63:0] _result_T_2329 = $signed(_result_T_2326) + $signed(_result_T_444);
  wire [63:0] _result_T_2332 = $signed(_result_T_2329) + $signed(_result_T_445);
  wire [63:0] _result_T_2335 = $signed(_result_T_2332) + $signed(_result_T_446);
  wire [63:0] _result_T_2338 = $signed(_result_T_2335) + $signed(_result_T_447);
  wire [63:0] _result_T_2341 = $signed(_result_T_2338) + $signed(_result_T_448);
  wire [63:0] _result_T_2344 = $signed(_result_T_2341) + $signed(_result_T_449);
  wire [63:0] _result_T_2347 = $signed(_result_T_2344) + $signed(_result_T_450);
  wire [63:0] _result_T_2350 = $signed(_result_T_2347) + $signed(_result_T_451);
  wire [63:0] _result_T_2353 = $signed(_result_T_2350) + $signed(_result_T_452);
  wire [63:0] _result_T_2356 = $signed(_result_T_2353) + $signed(_result_T_453);
  wire [63:0] _result_T_2359 = $signed(_result_T_2356) + $signed(_result_T_454);
  wire [63:0] _result_T_2362 = $signed(_result_T_2359) + $signed(_result_T_455);
  wire [63:0] _result_T_2365 = $signed(_result_T_2362) + $signed(_result_T_456);
  wire [63:0] _result_T_2368 = $signed(_result_T_2365) + $signed(_result_T_457);
  wire [63:0] _result_T_2371 = $signed(_result_T_2368) + $signed(_result_T_458);
  wire [63:0] _result_T_2374 = $signed(_result_T_2371) + $signed(_result_T_459);
  wire [63:0] _result_T_2377 = $signed(_result_T_2374) + $signed(_result_T_460);
  wire [63:0] _result_T_2380 = $signed(_result_T_2377) + $signed(_result_T_461);
  wire [63:0] _result_T_2383 = $signed(_result_T_2380) + $signed(_result_T_462);
  wire [63:0] _result_T_2386 = $signed(_result_T_2383) + $signed(_result_T_463);
  wire [63:0] _result_T_2389 = $signed(_result_T_2386) + $signed(_result_T_464);
  wire [63:0] _result_T_2392 = $signed(_result_T_2389) + $signed(_result_T_465);
  wire [63:0] _result_T_2395 = $signed(_result_T_2392) + $signed(_result_T_466);
  wire [63:0] _result_T_2398 = $signed(_result_T_2395) + $signed(_result_T_467);
  wire [63:0] _result_T_2401 = $signed(_result_T_2398) + $signed(_result_T_468);
  wire [63:0] _result_T_2404 = $signed(_result_T_2401) + $signed(_result_T_469);
  wire [63:0] _result_T_2407 = $signed(_result_T_2404) + $signed(_result_T_470);
  wire [63:0] _result_T_2410 = $signed(_result_T_2407) + $signed(_result_T_471);
  wire [63:0] _result_T_2413 = $signed(_result_T_2410) + $signed(_result_T_472);
  wire [63:0] _result_T_2416 = $signed(_result_T_2413) + $signed(_result_T_473);
  wire [63:0] _result_T_2419 = $signed(_result_T_2416) + $signed(_result_T_474);
  wire [63:0] _result_T_2422 = $signed(_result_T_2419) + $signed(_result_T_475);
  wire [63:0] _result_T_2425 = $signed(_result_T_2422) + $signed(_result_T_476);
  wire [63:0] _result_T_2428 = $signed(_result_T_2425) + $signed(_result_T_477);
  wire [63:0] _result_T_2431 = $signed(_result_T_2428) + $signed(_result_T_478);
  wire [63:0] _result_T_2434 = $signed(_result_T_2431) + $signed(_result_T_479);
  wire [63:0] _result_T_2437 = $signed(_result_T_2434) + $signed(_result_T_480);
  wire [63:0] _result_T_2440 = $signed(_result_T_2437) + $signed(_result_T_481);
  wire [63:0] _result_T_2443 = $signed(_result_T_2440) + $signed(_result_T_482);
  wire [63:0] _result_T_2446 = $signed(_result_T_2443) + $signed(_result_T_483);
  wire [63:0] _result_T_2449 = $signed(_result_T_2446) + $signed(_result_T_484);
  wire [63:0] _result_T_2452 = $signed(_result_T_2449) + $signed(_result_T_485);
  wire [63:0] _result_T_2455 = $signed(_result_T_2452) + $signed(_result_T_486);
  wire [63:0] _result_T_2458 = $signed(_result_T_2455) + $signed(_result_T_487);
  wire [63:0] _result_T_2461 = $signed(_result_T_2458) + $signed(_result_T_488);
  wire [63:0] _result_T_2464 = $signed(_result_T_2461) + $signed(_result_T_489);
  wire [63:0] _result_T_2467 = $signed(_result_T_2464) + $signed(_result_T_490);
  wire [63:0] _result_T_2470 = $signed(_result_T_2467) + $signed(_result_T_491);
  wire [63:0] _result_T_2473 = $signed(_result_T_2470) + $signed(_result_T_492);
  wire [63:0] _result_T_2476 = $signed(_result_T_2473) + $signed(_result_T_493);
  wire [63:0] _result_T_2479 = $signed(_result_T_2476) + $signed(_result_T_494);
  wire [63:0] _result_T_2482 = $signed(_result_T_2479) + $signed(_result_T_495);
  wire [63:0] _result_T_2485 = $signed(_result_T_2482) + $signed(_result_T_496);
  wire [63:0] _result_T_2488 = $signed(_result_T_2485) + $signed(_result_T_497);
  wire [63:0] _result_T_2491 = $signed(_result_T_2488) + $signed(_result_T_498);
  wire [63:0] _result_T_2494 = $signed(_result_T_2491) + $signed(_result_T_499);
  wire [63:0] _result_T_2497 = $signed(_result_T_2494) + $signed(_result_T_500);
  wire [63:0] _result_T_2500 = $signed(_result_T_2497) + $signed(_result_T_501);
  wire [63:0] _result_T_2503 = $signed(_result_T_2500) + $signed(_result_T_502);
  wire [63:0] _result_T_2506 = $signed(_result_T_2503) + $signed(_result_T_503);
  wire [63:0] _result_T_2509 = $signed(_result_T_2506) + $signed(_result_T_504);
  wire [63:0] _result_T_2512 = $signed(_result_T_2509) + $signed(_result_T_505);
  wire [63:0] _result_T_2515 = $signed(_result_T_2512) + $signed(_result_T_506);
  wire [63:0] _result_T_2518 = $signed(_result_T_2515) + $signed(_result_T_507);
  wire [63:0] _result_T_2521 = $signed(_result_T_2518) + $signed(_result_T_508);
  wire [63:0] _result_T_2524 = $signed(_result_T_2521) + $signed(_result_T_509);
  wire [63:0] _result_T_2527 = $signed(_result_T_2524) + $signed(_result_T_510);
  wire [63:0] _result_T_2530 = $signed(_result_T_2527) + $signed(_result_T_511);
  wire [63:0] _result_T_2533 = $signed(_result_T_2530) + $signed(_result_T_512);
  wire [63:0] _result_T_2536 = $signed(_result_T_2533) + $signed(_result_T_513);
  wire [63:0] _result_T_2539 = $signed(_result_T_2536) + $signed(_result_T_514);
  wire [63:0] _result_T_2542 = $signed(_result_T_2539) + $signed(_result_T_515);
  wire [63:0] _result_T_2545 = $signed(_result_T_2542) + $signed(_result_T_516);
  wire [63:0] _result_T_2548 = $signed(_result_T_2545) + $signed(_result_T_517);
  wire [63:0] _result_T_2551 = $signed(_result_T_2548) + $signed(_result_T_518);
  wire [63:0] _result_T_2554 = $signed(_result_T_2551) + $signed(_result_T_519);
  wire [63:0] _result_T_2557 = $signed(_result_T_2554) + $signed(_result_T_520);
  wire [63:0] _result_T_2560 = $signed(_result_T_2557) + $signed(_result_T_521);
  wire [63:0] _result_T_2563 = $signed(_result_T_2560) + $signed(_result_T_522);
  wire [63:0] _result_T_2566 = $signed(_result_T_2563) + $signed(_result_T_523);
  wire [63:0] _result_T_2569 = $signed(_result_T_2566) + $signed(_result_T_524);
  wire [63:0] _result_T_2572 = $signed(_result_T_2569) + $signed(_result_T_525);
  wire [63:0] _result_T_2575 = $signed(_result_T_2572) + $signed(_result_T_526);
  wire [63:0] _result_T_2578 = $signed(_result_T_2575) + $signed(_result_T_527);
  wire [63:0] _result_T_2581 = $signed(_result_T_2578) + $signed(_result_T_528);
  wire [63:0] _result_T_2584 = $signed(_result_T_2581) + $signed(_result_T_529);
  wire [63:0] _result_T_2587 = $signed(_result_T_2584) + $signed(_result_T_530);
  wire [63:0] _result_T_2590 = $signed(_result_T_2587) + $signed(_result_T_531);
  wire [63:0] _result_T_2593 = $signed(_result_T_2590) + $signed(_result_T_532);
  wire [63:0] _result_T_2596 = $signed(_result_T_2593) + $signed(_result_T_533);
  wire [63:0] _result_T_2599 = $signed(_result_T_2596) + $signed(_result_T_534);
  wire [63:0] _result_T_2602 = $signed(_result_T_2599) + $signed(_result_T_535);
  wire [63:0] _result_T_2605 = $signed(_result_T_2602) + $signed(_result_T_536);
  wire [63:0] _result_T_2608 = $signed(_result_T_2605) + $signed(_result_T_537);
  wire [63:0] _result_T_2611 = $signed(_result_T_2608) + $signed(_result_T_538);
  wire [63:0] _result_T_2614 = $signed(_result_T_2611) + $signed(_result_T_539);
  wire [63:0] _result_T_2617 = $signed(_result_T_2614) + $signed(_result_T_540);
  wire [63:0] _result_T_2620 = $signed(_result_T_2617) + $signed(_result_T_541);
  wire [63:0] _result_T_2623 = $signed(_result_T_2620) + $signed(_result_T_542);
  wire [63:0] _result_T_2626 = $signed(_result_T_2623) + $signed(_result_T_543);
  wire [63:0] _result_T_2629 = $signed(_result_T_2626) + $signed(_result_T_544);
  wire [63:0] _result_T_2632 = $signed(_result_T_2629) + $signed(_result_T_545);
  wire [63:0] _result_T_2635 = $signed(_result_T_2632) + $signed(_result_T_546);
  wire [63:0] _result_T_2638 = $signed(_result_T_2635) + $signed(_result_T_547);
  wire [63:0] _result_T_2641 = $signed(_result_T_2638) + $signed(_result_T_548);
  wire [63:0] _result_T_2644 = $signed(_result_T_2641) + $signed(_result_T_549);
  wire [63:0] _result_T_2647 = $signed(_result_T_2644) + $signed(_result_T_550);
  wire [63:0] _result_T_2650 = $signed(_result_T_2647) + $signed(_result_T_551);
  wire [63:0] _result_T_2653 = $signed(_result_T_2650) + $signed(_result_T_552);
  wire [63:0] _result_T_2656 = $signed(_result_T_2653) + $signed(_result_T_553);
  wire [63:0] _result_T_2659 = $signed(_result_T_2656) + $signed(_result_T_554);
  wire [63:0] _result_T_2662 = $signed(_result_T_2659) + $signed(_result_T_555);
  wire [63:0] _result_T_2665 = $signed(_result_T_2662) + $signed(_result_T_556);
  wire [63:0] _result_T_2668 = $signed(_result_T_2665) + $signed(_result_T_557);
  wire [63:0] _result_T_2671 = $signed(_result_T_2668) + $signed(_result_T_558);
  wire [63:0] _result_T_2674 = $signed(_result_T_2671) + $signed(_result_T_559);
  wire [63:0] _result_T_2677 = $signed(_result_T_2674) + $signed(_result_T_560);
  wire [63:0] _result_T_2680 = $signed(_result_T_2677) + $signed(_result_T_561);
  wire [63:0] _result_T_2683 = $signed(_result_T_2680) + $signed(_result_T_562);
  wire [63:0] _result_T_2686 = $signed(_result_T_2683) + $signed(_result_T_563);
  wire [63:0] _result_T_2689 = $signed(_result_T_2686) + $signed(_result_T_564);
  wire [63:0] _result_T_2692 = $signed(_result_T_2689) + $signed(_result_T_565);
  wire [63:0] _result_T_2695 = $signed(_result_T_2692) + $signed(_result_T_566);
  wire [63:0] _result_T_2698 = $signed(_result_T_2695) + $signed(_result_T_567);
  wire [63:0] _result_T_2701 = $signed(_result_T_2698) + $signed(_result_T_568);
  wire [63:0] _result_T_2704 = $signed(_result_T_2701) + $signed(_result_T_569);
  wire [63:0] _result_T_2707 = $signed(_result_T_2704) + $signed(_result_T_570);
  wire [63:0] _result_T_2710 = $signed(_result_T_2707) + $signed(_result_T_571);
  wire [63:0] _result_T_2713 = $signed(_result_T_2710) + $signed(_result_T_572);
  wire [63:0] _result_T_2716 = $signed(_result_T_2713) + $signed(_result_T_573);
  wire [63:0] _result_T_2719 = $signed(_result_T_2716) + $signed(_result_T_574);
  wire [63:0] _result_T_2722 = $signed(_result_T_2719) + $signed(_result_T_575);
  wire [63:0] _result_T_2725 = $signed(_result_T_2722) + $signed(_result_T_576);
  wire [63:0] _result_T_2728 = $signed(_result_T_2725) + $signed(_result_T_577);
  wire [63:0] _result_T_2731 = $signed(_result_T_2728) + $signed(_result_T_578);
  wire [63:0] _result_T_2734 = $signed(_result_T_2731) + $signed(_result_T_579);
  wire [63:0] _result_T_2737 = $signed(_result_T_2734) + $signed(_result_T_580);
  wire [63:0] _result_T_2740 = $signed(_result_T_2737) + $signed(_result_T_581);
  wire [63:0] _result_T_2743 = $signed(_result_T_2740) + $signed(_result_T_582);
  wire [63:0] _result_T_2746 = $signed(_result_T_2743) + $signed(_result_T_583);
  wire [63:0] _result_T_2749 = $signed(_result_T_2746) + $signed(_result_T_584);
  wire [63:0] _result_T_2752 = $signed(_result_T_2749) + $signed(_result_T_585);
  wire [63:0] _result_T_2755 = $signed(_result_T_2752) + $signed(_result_T_586);
  wire [63:0] _result_T_2758 = $signed(_result_T_2755) + $signed(_result_T_587);
  wire [63:0] _result_T_2761 = $signed(_result_T_2758) + $signed(_result_T_588);
  wire [63:0] _result_T_2764 = $signed(_result_T_2761) + $signed(_result_T_589);
  wire [63:0] _result_T_2767 = $signed(_result_T_2764) + $signed(_result_T_590);
  wire [63:0] _result_T_2770 = $signed(_result_T_2767) + $signed(_result_T_591);
  wire [63:0] _result_T_2773 = $signed(_result_T_2770) + $signed(_result_T_592);
  wire [63:0] _result_T_2776 = $signed(_result_T_2773) + $signed(_result_T_593);
  wire [63:0] _result_T_2779 = $signed(_result_T_2776) + $signed(_result_T_594);
  wire [63:0] _result_T_2782 = $signed(_result_T_2779) + $signed(_result_T_595);
  wire [63:0] _result_T_2785 = $signed(_result_T_2782) + $signed(_result_T_596);
  wire [63:0] _result_T_2788 = $signed(_result_T_2785) + $signed(_result_T_597);
  wire [63:0] _result_T_2791 = $signed(_result_T_2788) + $signed(_result_T_598);
  wire [63:0] _result_T_2794 = $signed(_result_T_2791) + $signed(_result_T_599);
  wire [63:0] _result_T_2797 = $signed(_result_T_2794) + $signed(_result_T_600);
  wire [63:0] _result_T_2800 = $signed(_result_T_2797) + $signed(_result_T_601);
  wire [63:0] _result_T_2803 = $signed(_result_T_2800) + $signed(_result_T_602);
  wire [63:0] _result_T_2806 = $signed(_result_T_2803) + $signed(_result_T_603);
  wire [63:0] _result_T_2809 = $signed(_result_T_2806) + $signed(_result_T_604);
  wire [63:0] _result_T_2812 = $signed(_result_T_2809) + $signed(_result_T_605);
  wire [63:0] _result_T_2815 = $signed(_result_T_2812) + $signed(_result_T_606);
  wire [63:0] _result_T_2818 = $signed(_result_T_2815) + $signed(_result_T_607);
  wire [63:0] _result_T_2821 = $signed(_result_T_2818) + $signed(_result_T_608);
  wire [63:0] _result_T_2824 = $signed(_result_T_2821) + $signed(_result_T_609);
  wire [63:0] _result_T_2827 = $signed(_result_T_2824) + $signed(_result_T_610);
  wire [63:0] _result_T_2830 = $signed(_result_T_2827) + $signed(_result_T_611);
  wire [63:0] _result_T_2833 = $signed(_result_T_2830) + $signed(_result_T_612);
  wire [63:0] _result_T_2836 = $signed(_result_T_2833) + $signed(_result_T_613);
  wire [63:0] _result_T_2839 = $signed(_result_T_2836) + $signed(_result_T_614);
  wire [63:0] _result_T_2842 = $signed(_result_T_2839) + $signed(_result_T_615);
  wire [63:0] _result_T_2845 = $signed(_result_T_2842) + $signed(_result_T_616);
  wire [63:0] _result_T_2848 = $signed(_result_T_2845) + $signed(_result_T_617);
  wire [63:0] _result_T_2851 = $signed(_result_T_2848) + $signed(_result_T_618);
  wire [63:0] _result_T_2854 = $signed(_result_T_2851) + $signed(_result_T_619);
  wire [63:0] _result_T_2857 = $signed(_result_T_2854) + $signed(_result_T_620);
  wire [63:0] _result_T_2860 = $signed(_result_T_2857) + $signed(_result_T_621);
  wire [63:0] _result_T_2863 = $signed(_result_T_2860) + $signed(_result_T_622);
  wire [63:0] _result_T_2866 = $signed(_result_T_2863) + $signed(_result_T_623);
  wire [63:0] _result_T_2869 = $signed(_result_T_2866) + $signed(_result_T_624);
  wire [63:0] _result_T_2872 = $signed(_result_T_2869) + $signed(_result_T_625);
  wire [63:0] _result_T_2875 = $signed(_result_T_2872) + $signed(_result_T_626);
  wire [63:0] _result_T_2878 = $signed(_result_T_2875) + $signed(_result_T_627);
  wire [63:0] _result_T_2881 = $signed(_result_T_2878) + $signed(_result_T_628);
  wire [63:0] _result_T_2884 = $signed(_result_T_2881) + $signed(_result_T_629);
  wire [63:0] _result_T_2887 = $signed(_result_T_2884) + $signed(_result_T_630);
  wire [63:0] _result_T_2890 = $signed(_result_T_2887) + $signed(_result_T_631);
  wire [63:0] _result_T_2893 = $signed(_result_T_2890) + $signed(_result_T_632);
  wire [63:0] _result_T_2896 = $signed(_result_T_2893) + $signed(_result_T_633);
  wire [63:0] _result_T_2899 = $signed(_result_T_2896) + $signed(_result_T_634);
  wire [63:0] _result_T_2902 = $signed(_result_T_2899) + $signed(_result_T_635);
  wire [63:0] _result_T_2905 = $signed(_result_T_2902) + $signed(_result_T_636);
  wire [63:0] _result_T_2908 = $signed(_result_T_2905) + $signed(_result_T_637);
  wire [63:0] _result_T_2911 = $signed(_result_T_2908) + $signed(_result_T_638);
  wire [63:0] _result_T_2914 = $signed(_result_T_2911) + $signed(_result_T_639);
  wire [63:0] _result_T_2917 = $signed(_result_T_2914) + $signed(_result_T_640);
  wire [63:0] _result_T_2920 = $signed(_result_T_2917) + $signed(_result_T_641);
  wire [63:0] _result_T_2923 = $signed(_result_T_2920) + $signed(_result_T_642);
  wire [63:0] _result_T_2926 = $signed(_result_T_2923) + $signed(_result_T_643);
  wire [63:0] _result_T_2929 = $signed(_result_T_2926) + $signed(_result_T_644);
  wire [63:0] _result_T_2932 = $signed(_result_T_2929) + $signed(_result_T_645);
  wire [63:0] _result_T_2935 = $signed(_result_T_2932) + $signed(_result_T_646);
  wire [63:0] _result_T_2938 = $signed(_result_T_2935) + $signed(_result_T_647);
  wire [63:0] _result_T_2941 = $signed(_result_T_2938) + $signed(_result_T_648);
  wire [63:0] _result_T_2944 = $signed(_result_T_2941) + $signed(_result_T_649);
  wire [63:0] _result_T_2947 = $signed(_result_T_2944) + $signed(_result_T_650);
  wire [63:0] _result_T_2950 = $signed(_result_T_2947) + $signed(_result_T_651);
  wire [63:0] _result_T_2953 = $signed(_result_T_2950) + $signed(_result_T_652);
  wire [63:0] _result_T_2956 = $signed(_result_T_2953) + $signed(_result_T_653);
  wire [63:0] _result_T_2959 = $signed(_result_T_2956) + $signed(_result_T_654);
  wire [63:0] _result_T_2962 = $signed(_result_T_2959) + $signed(_result_T_655);
  wire [63:0] _result_T_2965 = $signed(_result_T_2962) + $signed(_result_T_656);
  wire [63:0] _result_T_2968 = $signed(_result_T_2965) + $signed(_result_T_657);
  wire [63:0] _result_T_2971 = $signed(_result_T_2968) + $signed(_result_T_658);
  wire [63:0] _result_T_2974 = $signed(_result_T_2971) + $signed(_result_T_659);
  wire [63:0] _result_T_2977 = $signed(_result_T_2974) + $signed(_result_T_660);
  wire [63:0] _result_T_2980 = $signed(_result_T_2977) + $signed(_result_T_661);
  wire [63:0] _result_T_2983 = $signed(_result_T_2980) + $signed(_result_T_662);
  wire [63:0] _result_T_2986 = $signed(_result_T_2983) + $signed(_result_T_663);
  wire [63:0] _result_T_2989 = $signed(_result_T_2986) + $signed(_result_T_664);
  wire [63:0] _result_T_2992 = $signed(_result_T_2989) + $signed(_result_T_665);
  wire [63:0] _result_T_2995 = $signed(_result_T_2992) + $signed(_result_T_666);
  wire [63:0] _result_T_2998 = $signed(_result_T_2995) + $signed(_result_T_667);
  wire [63:0] _result_T_3001 = $signed(_result_T_2998) + $signed(_result_T_668);
  wire [63:0] _result_T_3004 = $signed(_result_T_3001) + $signed(_result_T_669);
  wire [63:0] _result_T_3007 = $signed(_result_T_3004) + $signed(_result_T_670);
  wire [63:0] _result_T_3010 = $signed(_result_T_3007) + $signed(_result_T_671);
  wire [63:0] _result_T_3013 = $signed(_result_T_3010) + $signed(_result_T_672);
  wire [63:0] _result_T_3016 = $signed(_result_T_3013) + $signed(_result_T_673);
  wire [63:0] _result_T_3019 = $signed(_result_T_3016) + $signed(_result_T_674);
  wire [63:0] _result_T_3022 = $signed(_result_T_3019) + $signed(_result_T_675);
  wire [63:0] _result_T_3025 = $signed(_result_T_3022) + $signed(_result_T_676);
  wire [63:0] _result_T_3028 = $signed(_result_T_3025) + $signed(_result_T_677);
  wire [63:0] _result_T_3031 = $signed(_result_T_3028) + $signed(_result_T_678);
  wire [63:0] _result_T_3034 = $signed(_result_T_3031) + $signed(_result_T_679);
  wire [63:0] _result_T_3037 = $signed(_result_T_3034) + $signed(_result_T_680);
  wire [63:0] _result_T_3040 = $signed(_result_T_3037) + $signed(_result_T_681);
  wire [63:0] _result_T_3043 = $signed(_result_T_3040) + $signed(_result_T_682);
  wire [63:0] _result_T_3046 = $signed(_result_T_3043) + $signed(_result_T_683);
  wire [63:0] _result_T_3049 = $signed(_result_T_3046) + $signed(_result_T_684);
  wire [63:0] _result_T_3052 = $signed(_result_T_3049) + $signed(_result_T_685);
  wire [63:0] _result_T_3055 = $signed(_result_T_3052) + $signed(_result_T_686);
  wire [63:0] _result_T_3058 = $signed(_result_T_3055) + $signed(_result_T_687);
  wire [63:0] _result_T_3061 = $signed(_result_T_3058) + $signed(_result_T_688);
  wire [63:0] _result_T_3064 = $signed(_result_T_3061) + $signed(_result_T_689);
  wire [63:0] _result_T_3067 = $signed(_result_T_3064) + $signed(_result_T_690);
  wire [63:0] _result_T_3070 = $signed(_result_T_3067) + $signed(_result_T_691);
  wire [63:0] _result_T_3073 = $signed(_result_T_3070) + $signed(_result_T_692);
  wire [63:0] _result_T_3076 = $signed(_result_T_3073) + $signed(_result_T_693);
  wire [63:0] _result_T_3079 = $signed(_result_T_3076) + $signed(_result_T_694);
  wire [63:0] _result_T_3082 = $signed(_result_T_3079) + $signed(_result_T_695);
  wire [63:0] _result_T_3085 = $signed(_result_T_3082) + $signed(_result_T_696);
  wire [63:0] _result_T_3088 = $signed(_result_T_3085) + $signed(_result_T_697);
  wire [63:0] _result_T_3091 = $signed(_result_T_3088) + $signed(_result_T_698);
  wire [63:0] _result_T_3094 = $signed(_result_T_3091) + $signed(_result_T_699);
  wire [63:0] _result_T_3097 = $signed(_result_T_3094) + $signed(_result_T_700);
  wire [63:0] _result_T_3100 = $signed(_result_T_3097) + $signed(_result_T_701);
  wire [63:0] _result_T_3103 = $signed(_result_T_3100) + $signed(_result_T_702);
  wire [63:0] _result_T_3106 = $signed(_result_T_3103) + $signed(_result_T_703);
  wire [63:0] _result_T_3109 = $signed(_result_T_3106) + $signed(_result_T_704);
  wire [63:0] _result_T_3112 = $signed(_result_T_3109) + $signed(_result_T_705);
  wire [63:0] _result_T_3115 = $signed(_result_T_3112) + $signed(_result_T_706);
  wire [63:0] _result_T_3118 = $signed(_result_T_3115) + $signed(_result_T_707);
  wire [63:0] _result_T_3121 = $signed(_result_T_3118) + $signed(_result_T_708);
  wire [63:0] _result_T_3124 = $signed(_result_T_3121) + $signed(_result_T_709);
  wire [63:0] _result_T_3127 = $signed(_result_T_3124) + $signed(_result_T_710);
  wire [63:0] _result_T_3130 = $signed(_result_T_3127) + $signed(_result_T_711);
  wire [63:0] _result_T_3133 = $signed(_result_T_3130) + $signed(_result_T_712);
  wire [63:0] _result_T_3136 = $signed(_result_T_3133) + $signed(_result_T_713);
  wire [63:0] _result_T_3139 = $signed(_result_T_3136) + $signed(_result_T_714);
  wire [63:0] _result_T_3142 = $signed(_result_T_3139) + $signed(_result_T_715);
  wire [63:0] _result_T_3145 = $signed(_result_T_3142) + $signed(_result_T_716);
  wire [63:0] _result_T_3148 = $signed(_result_T_3145) + $signed(_result_T_717);
  wire [63:0] _result_T_3151 = $signed(_result_T_3148) + $signed(_result_T_718);
  wire [63:0] _result_T_3154 = $signed(_result_T_3151) + $signed(_result_T_719);
  wire [63:0] _result_T_3157 = $signed(_result_T_3154) + $signed(_result_T_720);
  wire [63:0] _result_T_3160 = $signed(_result_T_3157) + $signed(_result_T_721);
  wire [63:0] _result_T_3163 = $signed(_result_T_3160) + $signed(_result_T_722);
  wire [63:0] _result_T_3166 = $signed(_result_T_3163) + $signed(_result_T_723);
  wire [63:0] _result_T_3169 = $signed(_result_T_3166) + $signed(_result_T_724);
  wire [63:0] _result_T_3172 = $signed(_result_T_3169) + $signed(_result_T_725);
  wire [63:0] _result_T_3175 = $signed(_result_T_3172) + $signed(_result_T_726);
  wire [63:0] _result_T_3178 = $signed(_result_T_3175) + $signed(_result_T_727);
  wire [63:0] _result_T_3181 = $signed(_result_T_3178) + $signed(_result_T_728);
  wire [63:0] _result_T_3184 = $signed(_result_T_3181) + $signed(_result_T_729);
  wire [63:0] _result_T_3187 = $signed(_result_T_3184) + $signed(_result_T_730);
  wire [63:0] _result_T_3190 = $signed(_result_T_3187) + $signed(_result_T_731);
  wire [63:0] _result_T_3193 = $signed(_result_T_3190) + $signed(_result_T_732);
  wire [63:0] _result_T_3196 = $signed(_result_T_3193) + $signed(_result_T_733);
  wire [63:0] _result_T_3199 = $signed(_result_T_3196) + $signed(_result_T_734);
  wire [63:0] _result_T_3202 = $signed(_result_T_3199) + $signed(_result_T_735);
  wire [63:0] _result_T_3205 = $signed(_result_T_3202) + $signed(_result_T_736);
  wire [63:0] _result_T_3208 = $signed(_result_T_3205) + $signed(_result_T_737);
  wire [63:0] _result_T_3211 = $signed(_result_T_3208) + $signed(_result_T_738);
  wire [63:0] _result_T_3214 = $signed(_result_T_3211) + $signed(_result_T_739);
  wire [63:0] _result_T_3217 = $signed(_result_T_3214) + $signed(_result_T_740);
  wire [63:0] _result_T_3220 = $signed(_result_T_3217) + $signed(_result_T_741);
  wire [63:0] _result_T_3223 = $signed(_result_T_3220) + $signed(_result_T_742);
  wire [63:0] _result_T_3226 = $signed(_result_T_3223) + $signed(_result_T_743);
  wire [63:0] _result_T_3229 = $signed(_result_T_3226) + $signed(_result_T_744);
  wire [63:0] _result_T_3232 = $signed(_result_T_3229) + $signed(_result_T_745);
  wire [63:0] _result_T_3235 = $signed(_result_T_3232) + $signed(_result_T_746);
  wire [63:0] _result_T_3238 = $signed(_result_T_3235) + $signed(_result_T_747);
  wire [63:0] _result_T_3241 = $signed(_result_T_3238) + $signed(_result_T_748);
  wire [63:0] _result_T_3244 = $signed(_result_T_3241) + $signed(_result_T_749);
  wire [63:0] _result_T_3247 = $signed(_result_T_3244) + $signed(_result_T_750);
  wire [63:0] _result_T_3250 = $signed(_result_T_3247) + $signed(_result_T_751);
  wire [63:0] _result_T_3253 = $signed(_result_T_3250) + $signed(_result_T_752);
  wire [63:0] _result_T_3256 = $signed(_result_T_3253) + $signed(_result_T_753);
  wire [63:0] _result_T_3259 = $signed(_result_T_3256) + $signed(_result_T_754);
  wire [63:0] _result_T_3262 = $signed(_result_T_3259) + $signed(_result_T_755);
  wire [63:0] _result_T_3265 = $signed(_result_T_3262) + $signed(_result_T_756);
  wire [63:0] _result_T_3268 = $signed(_result_T_3265) + $signed(_result_T_757);
  wire [63:0] _result_T_3271 = $signed(_result_T_3268) + $signed(_result_T_758);
  wire [63:0] _result_T_3274 = $signed(_result_T_3271) + $signed(_result_T_759);
  wire [63:0] _result_T_3277 = $signed(_result_T_3274) + $signed(_result_T_760);
  wire [63:0] _result_T_3280 = $signed(_result_T_3277) + $signed(_result_T_761);
  wire [63:0] _result_T_3283 = $signed(_result_T_3280) + $signed(_result_T_762);
  wire [63:0] _result_T_3286 = $signed(_result_T_3283) + $signed(_result_T_763);
  wire [63:0] _result_T_3289 = $signed(_result_T_3286) + $signed(_result_T_764);
  wire [63:0] _result_T_3292 = $signed(_result_T_3289) + $signed(_result_T_765);
  wire [63:0] _result_T_3295 = $signed(_result_T_3292) + $signed(_result_T_766);
  wire [63:0] _result_T_3298 = $signed(_result_T_3295) + $signed(_result_T_767);
  wire [63:0] _result_T_3301 = $signed(_result_T_3298) + $signed(_result_T_768);
  wire [63:0] _result_T_3304 = $signed(_result_T_3301) + $signed(_result_T_769);
  wire [63:0] _result_T_3307 = $signed(_result_T_3304) + $signed(_result_T_770);
  wire [63:0] _result_T_3310 = $signed(_result_T_3307) + $signed(_result_T_771);
  wire [63:0] _result_T_3313 = $signed(_result_T_3310) + $signed(_result_T_772);
  wire [63:0] _result_T_3316 = $signed(_result_T_3313) + $signed(_result_T_773);
  wire [63:0] _result_T_3319 = $signed(_result_T_3316) + $signed(_result_T_774);
  wire [63:0] _result_T_3322 = $signed(_result_T_3319) + $signed(_result_T_775);
  wire [63:0] _result_T_3325 = $signed(_result_T_3322) + $signed(_result_T_776);
  wire [63:0] _result_T_3328 = $signed(_result_T_3325) + $signed(_result_T_777);
  wire [63:0] _result_T_3331 = $signed(_result_T_3328) + $signed(_result_T_778);
  wire [63:0] _result_T_3334 = $signed(_result_T_3331) + $signed(_result_T_779);
  wire [63:0] _result_T_3337 = $signed(_result_T_3334) + $signed(_result_T_780);
  wire [63:0] _result_T_3340 = $signed(_result_T_3337) + $signed(_result_T_781);
  wire [63:0] _result_T_3343 = $signed(_result_T_3340) + $signed(_result_T_782);
  wire [63:0] _result_T_3346 = $signed(_result_T_3343) + $signed(_result_T_783);
  wire [63:0] _result_T_3349 = $signed(_result_T_3346) + $signed(_result_T_784);
  wire [63:0] _result_T_3352 = $signed(_result_T_3349) + $signed(_result_T_785);
  wire [63:0] _result_T_3355 = $signed(_result_T_3352) + $signed(_result_T_786);
  wire [63:0] _result_T_3358 = $signed(_result_T_3355) + $signed(_result_T_787);
  wire [63:0] _result_T_3361 = $signed(_result_T_3358) + $signed(_result_T_788);
  wire [63:0] _result_T_3364 = $signed(_result_T_3361) + $signed(_result_T_789);
  wire [63:0] _result_T_3367 = $signed(_result_T_3364) + $signed(_result_T_790);
  wire [63:0] _result_T_3370 = $signed(_result_T_3367) + $signed(_result_T_791);
  wire [63:0] _result_T_3373 = $signed(_result_T_3370) + $signed(_result_T_792);
  wire [63:0] _result_T_3376 = $signed(_result_T_3373) + $signed(_result_T_793);
  wire [63:0] _result_T_3379 = $signed(_result_T_3376) + $signed(_result_T_794);
  wire [63:0] _result_T_3382 = $signed(_result_T_3379) + $signed(_result_T_795);
  wire [63:0] _result_T_3385 = $signed(_result_T_3382) + $signed(_result_T_796);
  wire [63:0] _result_T_3388 = $signed(_result_T_3385) + $signed(_result_T_797);
  wire [63:0] _result_T_3391 = $signed(_result_T_3388) + $signed(_result_T_798);
  wire [63:0] _result_T_3394 = $signed(_result_T_3391) + $signed(_result_T_799);
  wire [63:0] _result_T_3397 = $signed(_result_T_3394) + $signed(_result_T_800);
  wire [63:0] _result_T_3400 = $signed(_result_T_3397) + $signed(_result_T_801);
  wire [63:0] _result_T_3403 = $signed(_result_T_3400) + $signed(_result_T_802);
  wire [63:0] _result_T_3406 = $signed(_result_T_3403) + $signed(_result_T_803);
  wire [63:0] _result_T_3409 = $signed(_result_T_3406) + $signed(_result_T_804);
  wire [63:0] _result_T_3412 = $signed(_result_T_3409) + $signed(_result_T_805);
  wire [63:0] _result_T_3415 = $signed(_result_T_3412) + $signed(_result_T_806);
  wire [63:0] _result_T_3418 = $signed(_result_T_3415) + $signed(_result_T_807);
  wire [63:0] _result_T_3421 = $signed(_result_T_3418) + $signed(_result_T_808);
  wire [63:0] _result_T_3424 = $signed(_result_T_3421) + $signed(_result_T_809);
  wire [63:0] _result_T_3427 = $signed(_result_T_3424) + $signed(_result_T_810);
  wire [63:0] _result_T_3430 = $signed(_result_T_3427) + $signed(_result_T_811);
  wire [63:0] _result_T_3433 = $signed(_result_T_3430) + $signed(_result_T_812);
  wire [63:0] _result_T_3436 = $signed(_result_T_3433) + $signed(_result_T_813);
  wire [63:0] _result_T_3439 = $signed(_result_T_3436) + $signed(_result_T_814);
  wire [63:0] _result_T_3442 = $signed(_result_T_3439) + $signed(_result_T_815);
  wire [63:0] _result_T_3445 = $signed(_result_T_3442) + $signed(_result_T_816);
  wire [63:0] _result_T_3448 = $signed(_result_T_3445) + $signed(_result_T_817);
  wire [63:0] _result_T_3451 = $signed(_result_T_3448) + $signed(_result_T_818);
  wire [63:0] _result_T_3454 = $signed(_result_T_3451) + $signed(_result_T_819);
  wire [63:0] _result_T_3457 = $signed(_result_T_3454) + $signed(_result_T_820);
  wire [63:0] _result_T_3460 = $signed(_result_T_3457) + $signed(_result_T_821);
  wire [63:0] _result_T_3463 = $signed(_result_T_3460) + $signed(_result_T_822);
  wire [63:0] _result_T_3466 = $signed(_result_T_3463) + $signed(_result_T_823);
  wire [63:0] _result_T_3469 = $signed(_result_T_3466) + $signed(_result_T_824);
  wire [63:0] _result_T_3472 = $signed(_result_T_3469) + $signed(_result_T_825);
  wire [63:0] _result_T_3475 = $signed(_result_T_3472) + $signed(_result_T_826);
  wire [63:0] _result_T_3478 = $signed(_result_T_3475) + $signed(_result_T_827);
  wire [63:0] _result_T_3481 = $signed(_result_T_3478) + $signed(_result_T_828);
  wire [63:0] _result_T_3484 = $signed(_result_T_3481) + $signed(_result_T_829);
  wire [63:0] _result_T_3487 = $signed(_result_T_3484) + $signed(_result_T_830);
  wire [63:0] _result_T_3490 = $signed(_result_T_3487) + $signed(_result_T_831);
  wire [63:0] _result_T_3493 = $signed(_result_T_3490) + $signed(_result_T_832);
  wire [63:0] _result_T_3496 = $signed(_result_T_3493) + $signed(_result_T_833);
  wire [63:0] _result_T_3499 = $signed(_result_T_3496) + $signed(_result_T_834);
  wire [63:0] _result_T_3502 = $signed(_result_T_3499) + $signed(_result_T_835);
  wire [63:0] _result_T_3505 = $signed(_result_T_3502) + $signed(_result_T_836);
  wire [63:0] _result_T_3508 = $signed(_result_T_3505) + $signed(_result_T_837);
  wire [63:0] _result_T_3511 = $signed(_result_T_3508) + $signed(_result_T_838);
  wire [63:0] _result_T_3514 = $signed(_result_T_3511) + $signed(_result_T_839);
  wire [63:0] _result_T_3517 = $signed(_result_T_3514) + $signed(_result_T_840);
  wire [63:0] _result_T_3520 = $signed(_result_T_3517) + $signed(_result_T_841);
  wire [63:0] _result_T_3523 = $signed(_result_T_3520) + $signed(_result_T_842);
  wire [63:0] _result_T_3526 = $signed(_result_T_3523) + $signed(_result_T_843);
  wire [63:0] _result_T_3529 = $signed(_result_T_3526) + $signed(_result_T_844);
  wire [63:0] _result_T_3532 = $signed(_result_T_3529) + $signed(_result_T_845);
  wire [63:0] _result_T_3535 = $signed(_result_T_3532) + $signed(_result_T_846);
  wire [63:0] _result_T_3538 = $signed(_result_T_3535) + $signed(_result_T_847);
  wire [63:0] _result_T_3541 = $signed(_result_T_3538) + $signed(_result_T_848);
  wire [63:0] _result_T_3544 = $signed(_result_T_3541) + $signed(_result_T_849);
  wire [63:0] _result_T_3547 = $signed(_result_T_3544) + $signed(_result_T_850);
  wire [63:0] _result_T_3550 = $signed(_result_T_3547) + $signed(_result_T_851);
  wire [63:0] _result_T_3553 = $signed(_result_T_3550) + $signed(_result_T_852);
  wire [63:0] _result_T_3556 = $signed(_result_T_3553) + $signed(_result_T_853);
  wire [63:0] _result_T_3559 = $signed(_result_T_3556) + $signed(_result_T_854);
  wire [63:0] _result_T_3562 = $signed(_result_T_3559) + $signed(_result_T_855);
  wire [63:0] _result_T_3565 = $signed(_result_T_3562) + $signed(_result_T_856);
  wire [63:0] _result_T_3568 = $signed(_result_T_3565) + $signed(_result_T_857);
  wire [63:0] _result_T_3571 = $signed(_result_T_3568) + $signed(_result_T_858);
  wire [63:0] _result_T_3574 = $signed(_result_T_3571) + $signed(_result_T_859);
  wire [63:0] _result_T_3577 = $signed(_result_T_3574) + $signed(_result_T_860);
  wire [63:0] _result_T_3580 = $signed(_result_T_3577) + $signed(_result_T_861);
  wire [63:0] _result_T_3583 = $signed(_result_T_3580) + $signed(_result_T_862);
  wire [63:0] _result_T_3586 = $signed(_result_T_3583) + $signed(_result_T_863);
  wire [63:0] _result_T_3589 = $signed(_result_T_3586) + $signed(_result_T_864);
  wire [63:0] _result_T_3592 = $signed(_result_T_3589) + $signed(_result_T_865);
  wire [63:0] _result_T_3595 = $signed(_result_T_3592) + $signed(_result_T_866);
  wire [63:0] _result_T_3598 = $signed(_result_T_3595) + $signed(_result_T_867);
  wire [63:0] _result_T_3601 = $signed(_result_T_3598) + $signed(_result_T_868);
  wire [63:0] _result_T_3604 = $signed(_result_T_3601) + $signed(_result_T_869);
  wire [63:0] _result_T_3607 = $signed(_result_T_3604) + $signed(_result_T_870);
  wire [63:0] _result_T_3610 = $signed(_result_T_3607) + $signed(_result_T_871);
  wire [63:0] _result_T_3613 = $signed(_result_T_3610) + $signed(_result_T_872);
  wire [63:0] _result_T_3616 = $signed(_result_T_3613) + $signed(_result_T_873);
  wire [63:0] _result_T_3619 = $signed(_result_T_3616) + $signed(_result_T_874);
  wire [63:0] _result_T_3622 = $signed(_result_T_3619) + $signed(_result_T_875);
  wire [63:0] _result_T_3625 = $signed(_result_T_3622) + $signed(_result_T_876);
  wire [63:0] _result_T_3628 = $signed(_result_T_3625) + $signed(_result_T_877);
  wire [63:0] _result_T_3631 = $signed(_result_T_3628) + $signed(_result_T_878);
  wire [63:0] _result_T_3634 = $signed(_result_T_3631) + $signed(_result_T_879);
  wire [63:0] _result_T_3637 = $signed(_result_T_3634) + $signed(_result_T_880);
  wire [63:0] _result_T_3640 = $signed(_result_T_3637) + $signed(_result_T_881);
  wire [63:0] _result_T_3643 = $signed(_result_T_3640) + $signed(_result_T_882);
  wire [63:0] _result_T_3646 = $signed(_result_T_3643) + $signed(_result_T_883);
  wire [63:0] _result_T_3649 = $signed(_result_T_3646) + $signed(_result_T_884);
  wire [63:0] _result_T_3652 = $signed(_result_T_3649) + $signed(_result_T_885);
  wire [63:0] _result_T_3655 = $signed(_result_T_3652) + $signed(_result_T_886);
  wire [63:0] _result_T_3658 = $signed(_result_T_3655) + $signed(_result_T_887);
  wire [63:0] _result_T_3661 = $signed(_result_T_3658) + $signed(_result_T_888);
  wire [63:0] _result_T_3664 = $signed(_result_T_3661) + $signed(_result_T_889);
  wire [63:0] _result_T_3667 = $signed(_result_T_3664) + $signed(_result_T_890);
  wire [63:0] _result_T_3670 = $signed(_result_T_3667) + $signed(_result_T_891);
  wire [63:0] _result_T_3673 = $signed(_result_T_3670) + $signed(_result_T_892);
  wire [63:0] _result_T_3676 = $signed(_result_T_3673) + $signed(_result_T_893);
  wire [63:0] _result_T_3679 = $signed(_result_T_3676) + $signed(_result_T_894);
  wire [63:0] _result_T_3682 = $signed(_result_T_3679) + $signed(_result_T_895);
  wire [63:0] _result_T_3685 = $signed(_result_T_3682) + $signed(_result_T_896);
  wire [63:0] _result_T_3688 = $signed(_result_T_3685) + $signed(_result_T_897);
  wire [63:0] _result_T_3691 = $signed(_result_T_3688) + $signed(_result_T_898);
  wire [63:0] _result_T_3694 = $signed(_result_T_3691) + $signed(_result_T_899);
  wire [63:0] _result_T_3697 = $signed(_result_T_3694) + $signed(_result_T_900);
  wire [63:0] _result_T_3700 = $signed(_result_T_3697) + $signed(_result_T_901);
  wire [63:0] _result_T_3703 = $signed(_result_T_3700) + $signed(_result_T_902);
  wire [63:0] _result_T_3706 = $signed(_result_T_3703) + $signed(_result_T_903);
  wire [63:0] _result_T_3709 = $signed(_result_T_3706) + $signed(_result_T_904);
  wire [63:0] _result_T_3712 = $signed(_result_T_3709) + $signed(_result_T_905);
  wire [63:0] _result_T_3715 = $signed(_result_T_3712) + $signed(_result_T_906);
  wire [63:0] _result_T_3718 = $signed(_result_T_3715) + $signed(_result_T_907);
  wire [63:0] _result_T_3721 = $signed(_result_T_3718) + $signed(_result_T_908);
  wire [63:0] _result_T_3724 = $signed(_result_T_3721) + $signed(_result_T_909);
  wire [63:0] _result_T_3727 = $signed(_result_T_3724) + $signed(_result_T_910);
  wire [63:0] _result_T_3730 = $signed(_result_T_3727) + $signed(_result_T_911);
  wire [63:0] _result_T_3733 = $signed(_result_T_3730) + $signed(_result_T_912);
  wire [63:0] _result_T_3736 = $signed(_result_T_3733) + $signed(_result_T_913);
  wire [63:0] _result_T_3739 = $signed(_result_T_3736) + $signed(_result_T_914);
  wire [63:0] _result_T_3742 = $signed(_result_T_3739) + $signed(_result_T_915);
  wire [63:0] _result_T_3745 = $signed(_result_T_3742) + $signed(_result_T_916);
  wire [63:0] _result_T_3748 = $signed(_result_T_3745) + $signed(_result_T_917);
  wire [63:0] _result_T_3751 = $signed(_result_T_3748) + $signed(_result_T_918);
  wire [63:0] _result_T_3754 = $signed(_result_T_3751) + $signed(_result_T_919);
  wire [63:0] _result_T_3757 = $signed(_result_T_3754) + $signed(_result_T_920);
  wire [63:0] _result_T_3760 = $signed(_result_T_3757) + $signed(_result_T_921);
  wire [63:0] _result_T_3763 = $signed(_result_T_3760) + $signed(_result_T_922);
  wire [63:0] _result_T_3766 = $signed(_result_T_3763) + $signed(_result_T_923);
  wire [63:0] _result_T_3769 = $signed(_result_T_3766) + $signed(_result_T_924);
  wire [63:0] _result_T_3772 = $signed(_result_T_3769) + $signed(_result_T_925);
  wire [63:0] _result_T_3775 = $signed(_result_T_3772) + $signed(_result_T_926);
  wire [63:0] _result_T_3778 = $signed(_result_T_3775) + $signed(_result_T_927);
  wire [63:0] _result_T_3781 = $signed(_result_T_3778) + $signed(_result_T_928);
  wire [63:0] _result_T_3784 = $signed(_result_T_3781) + $signed(_result_T_929);
  wire [63:0] _result_T_3787 = $signed(_result_T_3784) + $signed(_result_T_930);
  wire [63:0] _result_T_3790 = $signed(_result_T_3787) + $signed(_result_T_931);
  wire [63:0] _result_T_3793 = $signed(_result_T_3790) + $signed(_result_T_932);
  wire [63:0] _result_T_3796 = $signed(_result_T_3793) + $signed(_result_T_933);
  wire [63:0] _result_T_3799 = $signed(_result_T_3796) + $signed(_result_T_934);
  wire [63:0] _result_T_3802 = $signed(_result_T_3799) + $signed(_result_T_935);
  wire [63:0] _result_T_3805 = $signed(_result_T_3802) + $signed(_result_T_936);
  wire [63:0] _result_T_3808 = $signed(_result_T_3805) + $signed(_result_T_937);
  wire [63:0] _result_T_3811 = $signed(_result_T_3808) + $signed(_result_T_938);
  wire [63:0] _result_T_3814 = $signed(_result_T_3811) + $signed(_result_T_939);
  wire [63:0] _result_T_3817 = $signed(_result_T_3814) + $signed(_result_T_940);
  wire [63:0] _result_T_3820 = $signed(_result_T_3817) + $signed(_result_T_941);
  wire [63:0] _result_T_3823 = $signed(_result_T_3820) + $signed(_result_T_942);
  wire [63:0] _result_T_3826 = $signed(_result_T_3823) + $signed(_result_T_943);
  wire [63:0] _result_T_3829 = $signed(_result_T_3826) + $signed(_result_T_944);
  wire [63:0] _result_T_3832 = $signed(_result_T_3829) + $signed(_result_T_945);
  wire [63:0] _result_T_3835 = $signed(_result_T_3832) + $signed(_result_T_946);
  wire [63:0] _result_T_3838 = $signed(_result_T_3835) + $signed(_result_T_947);
  wire [63:0] _result_T_3841 = $signed(_result_T_3838) + $signed(_result_T_948);
  wire [63:0] _result_T_3844 = $signed(_result_T_3841) + $signed(_result_T_949);
  wire [63:0] _result_T_3847 = $signed(_result_T_3844) + $signed(_result_T_950);
  wire [63:0] _result_T_3850 = $signed(_result_T_3847) + $signed(_result_T_951);
  wire [63:0] _result_T_3853 = $signed(_result_T_3850) + $signed(_result_T_952);
  wire [63:0] _result_T_3856 = $signed(_result_T_3853) + $signed(_result_T_953);
  wire [63:0] _result_T_3859 = $signed(_result_T_3856) + $signed(_result_T_954);
  wire [63:0] _result_T_3862 = $signed(_result_T_3859) + $signed(_result_T_955);
  wire [63:0] _result_T_3865 = $signed(_result_T_3862) + $signed(_result_T_956);
  wire [63:0] _result_T_3868 = $signed(_result_T_3865) + $signed(_result_T_957);
  wire [63:0] _result_T_3871 = $signed(_result_T_3868) + $signed(_result_T_958);
  wire [63:0] _result_T_3874 = $signed(_result_T_3871) + $signed(_result_T_959);
  wire [63:0] _result_T_3877 = $signed(_result_T_3874) + $signed(_result_T_960);
  wire [63:0] _result_T_3880 = $signed(_result_T_3877) + $signed(_result_T_961);
  wire [63:0] _result_T_3883 = $signed(_result_T_3880) + $signed(_result_T_962);
  wire [63:0] _result_T_3886 = $signed(_result_T_3883) + $signed(_result_T_963);
  wire [63:0] _result_T_3889 = $signed(_result_T_3886) + $signed(_result_T_964);
  wire [63:0] _result_T_3892 = $signed(_result_T_3889) + $signed(_result_T_965);
  wire [63:0] _result_T_3895 = $signed(_result_T_3892) + $signed(_result_T_966);
  wire [63:0] _result_T_3898 = $signed(_result_T_3895) + $signed(_result_T_967);
  wire [63:0] _result_T_3901 = $signed(_result_T_3898) + $signed(_result_T_968);
  wire [63:0] _result_T_3904 = $signed(_result_T_3901) + $signed(_result_T_969);
  wire [63:0] _result_T_3907 = $signed(_result_T_3904) + $signed(_result_T_970);
  wire [63:0] _result_T_3910 = $signed(_result_T_3907) + $signed(_result_T_971);
  wire [63:0] _result_T_3913 = $signed(_result_T_3910) + $signed(_result_T_972);
  wire [63:0] _result_T_3916 = $signed(_result_T_3913) + $signed(_result_T_973);
  wire [63:0] _result_T_3919 = $signed(_result_T_3916) + $signed(_result_T_974);
  wire [63:0] _result_T_3922 = $signed(_result_T_3919) + $signed(_result_T_975);
  wire [63:0] _result_T_3925 = $signed(_result_T_3922) + $signed(_result_T_976);
  wire [63:0] _result_T_3928 = $signed(_result_T_3925) + $signed(_result_T_977);
  wire [63:0] _result_T_3931 = $signed(_result_T_3928) + $signed(_result_T_978);
  wire [63:0] _result_T_3934 = $signed(_result_T_3931) + $signed(_result_T_979);
  wire [63:0] _result_T_3937 = $signed(_result_T_3934) + $signed(_result_T_980);
  wire [63:0] _result_T_3940 = $signed(_result_T_3937) + $signed(_result_T_981);
  wire [63:0] _result_T_3943 = $signed(_result_T_3940) + $signed(_result_T_982);
  wire [63:0] _result_T_3946 = $signed(_result_T_3943) + $signed(_result_T_983);
  wire [63:0] _result_T_3949 = $signed(_result_T_3946) + $signed(_result_T_984);
  wire [63:0] _result_T_3952 = $signed(_result_T_3949) + $signed(_result_T_985);
  wire [63:0] _result_T_3955 = $signed(_result_T_3952) + $signed(_result_T_986);
  wire [63:0] _result_T_3958 = $signed(_result_T_3955) + $signed(_result_T_987);
  wire [63:0] _result_T_3961 = $signed(_result_T_3958) + $signed(_result_T_988);
  wire [63:0] _result_T_3964 = $signed(_result_T_3961) + $signed(_result_T_989);
  wire [63:0] _result_T_3967 = $signed(_result_T_3964) + $signed(_result_T_990);
  wire [63:0] _result_T_3970 = $signed(_result_T_3967) + $signed(_result_T_991);
  wire [63:0] _result_T_3973 = $signed(_result_T_3970) + $signed(_result_T_992);
  wire [63:0] _result_T_3976 = $signed(_result_T_3973) + $signed(_result_T_993);
  wire [63:0] _result_T_3979 = $signed(_result_T_3976) + $signed(_result_T_994);
  wire [63:0] _result_T_3982 = $signed(_result_T_3979) + $signed(_result_T_995);
  wire [63:0] _result_T_3985 = $signed(_result_T_3982) + $signed(_result_T_996);
  wire [63:0] _result_T_3988 = $signed(_result_T_3985) + $signed(_result_T_997);
  wire [63:0] _result_T_3991 = $signed(_result_T_3988) + $signed(_result_T_998);
  wire [63:0] _result_T_3994 = $signed(_result_T_3991) + $signed(_result_T_999);
  wire [63:0] _result_T_3997 = $signed(_result_T_3994) + $signed(_result_T_1000);
  wire [79:0] _GEN_1000 = insn[6:0] == 7'h5b ? $signed({{16{_result_T_3997[63]}},_result_T_3997}) : $signed({$signed(
    result), 16'h0});
  wire [79:0] _GEN_2001 = insn[6:0] == 7'h2b ? $signed({$signed(result), 16'h0}) : $signed(_GEN_1000);
  wire [79:0] _GEN_4002 = insn[6:0] == 7'hb ? $signed({$signed(result), 16'h0}) : $signed(_GEN_2001);
  wire [79:0] _GEN_6003 = valid ? $signed(_GEN_4002) : $signed({$signed(result), 16'h0});
  assign rd = result[31:0];
  always @(posedge clock) begin
    if (reset) begin
      coeffs_0 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h0 == rs2[9:0]) begin
          coeffs_0 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_1 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1 == rs2[9:0]) begin
          coeffs_1 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_2 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2 == rs2[9:0]) begin
          coeffs_2 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_3 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3 == rs2[9:0]) begin
          coeffs_3 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_4 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h4 == rs2[9:0]) begin
          coeffs_4 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_5 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h5 == rs2[9:0]) begin
          coeffs_5 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_6 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h6 == rs2[9:0]) begin
          coeffs_6 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_7 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h7 == rs2[9:0]) begin
          coeffs_7 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_8 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h8 == rs2[9:0]) begin
          coeffs_8 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_9 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h9 == rs2[9:0]) begin
          coeffs_9 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_10 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha == rs2[9:0]) begin
          coeffs_10 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_11 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb == rs2[9:0]) begin
          coeffs_11 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_12 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc == rs2[9:0]) begin
          coeffs_12 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_13 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd == rs2[9:0]) begin
          coeffs_13 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_14 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he == rs2[9:0]) begin
          coeffs_14 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_15 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf == rs2[9:0]) begin
          coeffs_15 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_16 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h10 == rs2[9:0]) begin
          coeffs_16 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_17 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h11 == rs2[9:0]) begin
          coeffs_17 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_18 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h12 == rs2[9:0]) begin
          coeffs_18 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_19 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h13 == rs2[9:0]) begin
          coeffs_19 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_20 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h14 == rs2[9:0]) begin
          coeffs_20 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_21 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h15 == rs2[9:0]) begin
          coeffs_21 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_22 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h16 == rs2[9:0]) begin
          coeffs_22 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_23 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h17 == rs2[9:0]) begin
          coeffs_23 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_24 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h18 == rs2[9:0]) begin
          coeffs_24 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_25 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h19 == rs2[9:0]) begin
          coeffs_25 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_26 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a == rs2[9:0]) begin
          coeffs_26 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_27 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b == rs2[9:0]) begin
          coeffs_27 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_28 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c == rs2[9:0]) begin
          coeffs_28 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_29 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d == rs2[9:0]) begin
          coeffs_29 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_30 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e == rs2[9:0]) begin
          coeffs_30 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_31 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f == rs2[9:0]) begin
          coeffs_31 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_32 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h20 == rs2[9:0]) begin
          coeffs_32 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_33 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h21 == rs2[9:0]) begin
          coeffs_33 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_34 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h22 == rs2[9:0]) begin
          coeffs_34 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_35 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h23 == rs2[9:0]) begin
          coeffs_35 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_36 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h24 == rs2[9:0]) begin
          coeffs_36 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_37 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h25 == rs2[9:0]) begin
          coeffs_37 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_38 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h26 == rs2[9:0]) begin
          coeffs_38 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_39 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h27 == rs2[9:0]) begin
          coeffs_39 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_40 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h28 == rs2[9:0]) begin
          coeffs_40 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_41 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h29 == rs2[9:0]) begin
          coeffs_41 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_42 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a == rs2[9:0]) begin
          coeffs_42 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_43 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b == rs2[9:0]) begin
          coeffs_43 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_44 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c == rs2[9:0]) begin
          coeffs_44 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_45 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d == rs2[9:0]) begin
          coeffs_45 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_46 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e == rs2[9:0]) begin
          coeffs_46 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_47 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f == rs2[9:0]) begin
          coeffs_47 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_48 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h30 == rs2[9:0]) begin
          coeffs_48 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_49 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h31 == rs2[9:0]) begin
          coeffs_49 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_50 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h32 == rs2[9:0]) begin
          coeffs_50 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_51 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h33 == rs2[9:0]) begin
          coeffs_51 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_52 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h34 == rs2[9:0]) begin
          coeffs_52 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_53 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h35 == rs2[9:0]) begin
          coeffs_53 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_54 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h36 == rs2[9:0]) begin
          coeffs_54 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_55 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h37 == rs2[9:0]) begin
          coeffs_55 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_56 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h38 == rs2[9:0]) begin
          coeffs_56 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_57 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h39 == rs2[9:0]) begin
          coeffs_57 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_58 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a == rs2[9:0]) begin
          coeffs_58 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_59 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b == rs2[9:0]) begin
          coeffs_59 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_60 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c == rs2[9:0]) begin
          coeffs_60 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_61 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d == rs2[9:0]) begin
          coeffs_61 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_62 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3e == rs2[9:0]) begin
          coeffs_62 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_63 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3f == rs2[9:0]) begin
          coeffs_63 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_64 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h40 == rs2[9:0]) begin
          coeffs_64 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_65 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h41 == rs2[9:0]) begin
          coeffs_65 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_66 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h42 == rs2[9:0]) begin
          coeffs_66 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_67 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h43 == rs2[9:0]) begin
          coeffs_67 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_68 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h44 == rs2[9:0]) begin
          coeffs_68 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_69 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h45 == rs2[9:0]) begin
          coeffs_69 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_70 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h46 == rs2[9:0]) begin
          coeffs_70 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_71 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h47 == rs2[9:0]) begin
          coeffs_71 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_72 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h48 == rs2[9:0]) begin
          coeffs_72 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_73 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h49 == rs2[9:0]) begin
          coeffs_73 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_74 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h4a == rs2[9:0]) begin
          coeffs_74 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_75 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h4b == rs2[9:0]) begin
          coeffs_75 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_76 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h4c == rs2[9:0]) begin
          coeffs_76 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_77 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h4d == rs2[9:0]) begin
          coeffs_77 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_78 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h4e == rs2[9:0]) begin
          coeffs_78 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_79 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h4f == rs2[9:0]) begin
          coeffs_79 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_80 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h50 == rs2[9:0]) begin
          coeffs_80 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_81 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h51 == rs2[9:0]) begin
          coeffs_81 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_82 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h52 == rs2[9:0]) begin
          coeffs_82 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_83 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h53 == rs2[9:0]) begin
          coeffs_83 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_84 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h54 == rs2[9:0]) begin
          coeffs_84 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_85 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h55 == rs2[9:0]) begin
          coeffs_85 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_86 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h56 == rs2[9:0]) begin
          coeffs_86 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_87 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h57 == rs2[9:0]) begin
          coeffs_87 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_88 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h58 == rs2[9:0]) begin
          coeffs_88 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_89 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h59 == rs2[9:0]) begin
          coeffs_89 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_90 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h5a == rs2[9:0]) begin
          coeffs_90 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_91 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h5b == rs2[9:0]) begin
          coeffs_91 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_92 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h5c == rs2[9:0]) begin
          coeffs_92 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_93 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h5d == rs2[9:0]) begin
          coeffs_93 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_94 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h5e == rs2[9:0]) begin
          coeffs_94 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_95 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h5f == rs2[9:0]) begin
          coeffs_95 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_96 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h60 == rs2[9:0]) begin
          coeffs_96 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_97 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h61 == rs2[9:0]) begin
          coeffs_97 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_98 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h62 == rs2[9:0]) begin
          coeffs_98 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_99 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h63 == rs2[9:0]) begin
          coeffs_99 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_100 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h64 == rs2[9:0]) begin
          coeffs_100 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_101 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h65 == rs2[9:0]) begin
          coeffs_101 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_102 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h66 == rs2[9:0]) begin
          coeffs_102 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_103 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h67 == rs2[9:0]) begin
          coeffs_103 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_104 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h68 == rs2[9:0]) begin
          coeffs_104 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_105 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h69 == rs2[9:0]) begin
          coeffs_105 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_106 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h6a == rs2[9:0]) begin
          coeffs_106 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_107 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h6b == rs2[9:0]) begin
          coeffs_107 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_108 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h6c == rs2[9:0]) begin
          coeffs_108 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_109 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h6d == rs2[9:0]) begin
          coeffs_109 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_110 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h6e == rs2[9:0]) begin
          coeffs_110 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_111 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h6f == rs2[9:0]) begin
          coeffs_111 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_112 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h70 == rs2[9:0]) begin
          coeffs_112 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_113 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h71 == rs2[9:0]) begin
          coeffs_113 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_114 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h72 == rs2[9:0]) begin
          coeffs_114 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_115 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h73 == rs2[9:0]) begin
          coeffs_115 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_116 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h74 == rs2[9:0]) begin
          coeffs_116 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_117 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h75 == rs2[9:0]) begin
          coeffs_117 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_118 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h76 == rs2[9:0]) begin
          coeffs_118 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_119 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h77 == rs2[9:0]) begin
          coeffs_119 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_120 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h78 == rs2[9:0]) begin
          coeffs_120 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_121 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h79 == rs2[9:0]) begin
          coeffs_121 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_122 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h7a == rs2[9:0]) begin
          coeffs_122 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_123 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h7b == rs2[9:0]) begin
          coeffs_123 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_124 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h7c == rs2[9:0]) begin
          coeffs_124 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_125 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h7d == rs2[9:0]) begin
          coeffs_125 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_126 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h7e == rs2[9:0]) begin
          coeffs_126 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_127 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h7f == rs2[9:0]) begin
          coeffs_127 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_128 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h80 == rs2[9:0]) begin
          coeffs_128 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_129 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h81 == rs2[9:0]) begin
          coeffs_129 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_130 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h82 == rs2[9:0]) begin
          coeffs_130 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_131 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h83 == rs2[9:0]) begin
          coeffs_131 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_132 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h84 == rs2[9:0]) begin
          coeffs_132 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_133 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h85 == rs2[9:0]) begin
          coeffs_133 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_134 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h86 == rs2[9:0]) begin
          coeffs_134 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_135 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h87 == rs2[9:0]) begin
          coeffs_135 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_136 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h88 == rs2[9:0]) begin
          coeffs_136 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_137 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h89 == rs2[9:0]) begin
          coeffs_137 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_138 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h8a == rs2[9:0]) begin
          coeffs_138 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_139 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h8b == rs2[9:0]) begin
          coeffs_139 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_140 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h8c == rs2[9:0]) begin
          coeffs_140 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_141 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h8d == rs2[9:0]) begin
          coeffs_141 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_142 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h8e == rs2[9:0]) begin
          coeffs_142 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_143 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h8f == rs2[9:0]) begin
          coeffs_143 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_144 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h90 == rs2[9:0]) begin
          coeffs_144 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_145 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h91 == rs2[9:0]) begin
          coeffs_145 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_146 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h92 == rs2[9:0]) begin
          coeffs_146 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_147 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h93 == rs2[9:0]) begin
          coeffs_147 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_148 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h94 == rs2[9:0]) begin
          coeffs_148 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_149 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h95 == rs2[9:0]) begin
          coeffs_149 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_150 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h96 == rs2[9:0]) begin
          coeffs_150 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_151 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h97 == rs2[9:0]) begin
          coeffs_151 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_152 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h98 == rs2[9:0]) begin
          coeffs_152 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_153 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h99 == rs2[9:0]) begin
          coeffs_153 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_154 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h9a == rs2[9:0]) begin
          coeffs_154 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_155 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h9b == rs2[9:0]) begin
          coeffs_155 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_156 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h9c == rs2[9:0]) begin
          coeffs_156 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_157 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h9d == rs2[9:0]) begin
          coeffs_157 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_158 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h9e == rs2[9:0]) begin
          coeffs_158 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_159 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h9f == rs2[9:0]) begin
          coeffs_159 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_160 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha0 == rs2[9:0]) begin
          coeffs_160 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_161 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha1 == rs2[9:0]) begin
          coeffs_161 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_162 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha2 == rs2[9:0]) begin
          coeffs_162 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_163 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha3 == rs2[9:0]) begin
          coeffs_163 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_164 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha4 == rs2[9:0]) begin
          coeffs_164 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_165 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha5 == rs2[9:0]) begin
          coeffs_165 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_166 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha6 == rs2[9:0]) begin
          coeffs_166 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_167 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha7 == rs2[9:0]) begin
          coeffs_167 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_168 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha8 == rs2[9:0]) begin
          coeffs_168 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_169 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha9 == rs2[9:0]) begin
          coeffs_169 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_170 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'haa == rs2[9:0]) begin
          coeffs_170 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_171 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hab == rs2[9:0]) begin
          coeffs_171 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_172 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hac == rs2[9:0]) begin
          coeffs_172 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_173 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'had == rs2[9:0]) begin
          coeffs_173 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_174 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hae == rs2[9:0]) begin
          coeffs_174 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_175 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'haf == rs2[9:0]) begin
          coeffs_175 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_176 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb0 == rs2[9:0]) begin
          coeffs_176 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_177 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb1 == rs2[9:0]) begin
          coeffs_177 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_178 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb2 == rs2[9:0]) begin
          coeffs_178 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_179 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb3 == rs2[9:0]) begin
          coeffs_179 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_180 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb4 == rs2[9:0]) begin
          coeffs_180 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_181 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb5 == rs2[9:0]) begin
          coeffs_181 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_182 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb6 == rs2[9:0]) begin
          coeffs_182 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_183 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb7 == rs2[9:0]) begin
          coeffs_183 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_184 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb8 == rs2[9:0]) begin
          coeffs_184 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_185 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb9 == rs2[9:0]) begin
          coeffs_185 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_186 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hba == rs2[9:0]) begin
          coeffs_186 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_187 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hbb == rs2[9:0]) begin
          coeffs_187 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_188 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hbc == rs2[9:0]) begin
          coeffs_188 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_189 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hbd == rs2[9:0]) begin
          coeffs_189 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_190 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hbe == rs2[9:0]) begin
          coeffs_190 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_191 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hbf == rs2[9:0]) begin
          coeffs_191 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_192 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc0 == rs2[9:0]) begin
          coeffs_192 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_193 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc1 == rs2[9:0]) begin
          coeffs_193 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_194 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc2 == rs2[9:0]) begin
          coeffs_194 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_195 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc3 == rs2[9:0]) begin
          coeffs_195 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_196 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc4 == rs2[9:0]) begin
          coeffs_196 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_197 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc5 == rs2[9:0]) begin
          coeffs_197 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_198 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc6 == rs2[9:0]) begin
          coeffs_198 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_199 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc7 == rs2[9:0]) begin
          coeffs_199 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_200 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc8 == rs2[9:0]) begin
          coeffs_200 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_201 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc9 == rs2[9:0]) begin
          coeffs_201 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_202 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hca == rs2[9:0]) begin
          coeffs_202 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_203 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hcb == rs2[9:0]) begin
          coeffs_203 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_204 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hcc == rs2[9:0]) begin
          coeffs_204 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_205 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hcd == rs2[9:0]) begin
          coeffs_205 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_206 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hce == rs2[9:0]) begin
          coeffs_206 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_207 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hcf == rs2[9:0]) begin
          coeffs_207 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_208 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd0 == rs2[9:0]) begin
          coeffs_208 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_209 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd1 == rs2[9:0]) begin
          coeffs_209 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_210 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd2 == rs2[9:0]) begin
          coeffs_210 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_211 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd3 == rs2[9:0]) begin
          coeffs_211 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_212 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd4 == rs2[9:0]) begin
          coeffs_212 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_213 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd5 == rs2[9:0]) begin
          coeffs_213 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_214 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd6 == rs2[9:0]) begin
          coeffs_214 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_215 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd7 == rs2[9:0]) begin
          coeffs_215 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_216 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd8 == rs2[9:0]) begin
          coeffs_216 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_217 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd9 == rs2[9:0]) begin
          coeffs_217 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_218 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hda == rs2[9:0]) begin
          coeffs_218 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_219 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hdb == rs2[9:0]) begin
          coeffs_219 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_220 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hdc == rs2[9:0]) begin
          coeffs_220 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_221 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hdd == rs2[9:0]) begin
          coeffs_221 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_222 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hde == rs2[9:0]) begin
          coeffs_222 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_223 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hdf == rs2[9:0]) begin
          coeffs_223 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_224 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he0 == rs2[9:0]) begin
          coeffs_224 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_225 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he1 == rs2[9:0]) begin
          coeffs_225 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_226 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he2 == rs2[9:0]) begin
          coeffs_226 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_227 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he3 == rs2[9:0]) begin
          coeffs_227 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_228 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he4 == rs2[9:0]) begin
          coeffs_228 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_229 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he5 == rs2[9:0]) begin
          coeffs_229 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_230 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he6 == rs2[9:0]) begin
          coeffs_230 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_231 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he7 == rs2[9:0]) begin
          coeffs_231 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_232 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he8 == rs2[9:0]) begin
          coeffs_232 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_233 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he9 == rs2[9:0]) begin
          coeffs_233 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_234 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hea == rs2[9:0]) begin
          coeffs_234 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_235 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'heb == rs2[9:0]) begin
          coeffs_235 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_236 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hec == rs2[9:0]) begin
          coeffs_236 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_237 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hed == rs2[9:0]) begin
          coeffs_237 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_238 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hee == rs2[9:0]) begin
          coeffs_238 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_239 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hef == rs2[9:0]) begin
          coeffs_239 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_240 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf0 == rs2[9:0]) begin
          coeffs_240 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_241 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf1 == rs2[9:0]) begin
          coeffs_241 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_242 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf2 == rs2[9:0]) begin
          coeffs_242 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_243 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf3 == rs2[9:0]) begin
          coeffs_243 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_244 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf4 == rs2[9:0]) begin
          coeffs_244 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_245 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf5 == rs2[9:0]) begin
          coeffs_245 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_246 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf6 == rs2[9:0]) begin
          coeffs_246 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_247 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf7 == rs2[9:0]) begin
          coeffs_247 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_248 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf8 == rs2[9:0]) begin
          coeffs_248 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_249 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf9 == rs2[9:0]) begin
          coeffs_249 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_250 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hfa == rs2[9:0]) begin
          coeffs_250 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_251 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hfb == rs2[9:0]) begin
          coeffs_251 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_252 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hfc == rs2[9:0]) begin
          coeffs_252 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_253 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hfd == rs2[9:0]) begin
          coeffs_253 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_254 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hfe == rs2[9:0]) begin
          coeffs_254 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_255 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hff == rs2[9:0]) begin
          coeffs_255 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_256 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h100 == rs2[9:0]) begin
          coeffs_256 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_257 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h101 == rs2[9:0]) begin
          coeffs_257 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_258 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h102 == rs2[9:0]) begin
          coeffs_258 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_259 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h103 == rs2[9:0]) begin
          coeffs_259 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_260 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h104 == rs2[9:0]) begin
          coeffs_260 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_261 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h105 == rs2[9:0]) begin
          coeffs_261 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_262 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h106 == rs2[9:0]) begin
          coeffs_262 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_263 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h107 == rs2[9:0]) begin
          coeffs_263 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_264 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h108 == rs2[9:0]) begin
          coeffs_264 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_265 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h109 == rs2[9:0]) begin
          coeffs_265 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_266 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h10a == rs2[9:0]) begin
          coeffs_266 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_267 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h10b == rs2[9:0]) begin
          coeffs_267 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_268 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h10c == rs2[9:0]) begin
          coeffs_268 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_269 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h10d == rs2[9:0]) begin
          coeffs_269 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_270 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h10e == rs2[9:0]) begin
          coeffs_270 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_271 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h10f == rs2[9:0]) begin
          coeffs_271 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_272 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h110 == rs2[9:0]) begin
          coeffs_272 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_273 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h111 == rs2[9:0]) begin
          coeffs_273 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_274 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h112 == rs2[9:0]) begin
          coeffs_274 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_275 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h113 == rs2[9:0]) begin
          coeffs_275 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_276 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h114 == rs2[9:0]) begin
          coeffs_276 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_277 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h115 == rs2[9:0]) begin
          coeffs_277 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_278 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h116 == rs2[9:0]) begin
          coeffs_278 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_279 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h117 == rs2[9:0]) begin
          coeffs_279 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_280 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h118 == rs2[9:0]) begin
          coeffs_280 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_281 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h119 == rs2[9:0]) begin
          coeffs_281 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_282 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h11a == rs2[9:0]) begin
          coeffs_282 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_283 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h11b == rs2[9:0]) begin
          coeffs_283 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_284 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h11c == rs2[9:0]) begin
          coeffs_284 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_285 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h11d == rs2[9:0]) begin
          coeffs_285 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_286 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h11e == rs2[9:0]) begin
          coeffs_286 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_287 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h11f == rs2[9:0]) begin
          coeffs_287 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_288 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h120 == rs2[9:0]) begin
          coeffs_288 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_289 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h121 == rs2[9:0]) begin
          coeffs_289 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_290 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h122 == rs2[9:0]) begin
          coeffs_290 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_291 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h123 == rs2[9:0]) begin
          coeffs_291 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_292 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h124 == rs2[9:0]) begin
          coeffs_292 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_293 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h125 == rs2[9:0]) begin
          coeffs_293 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_294 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h126 == rs2[9:0]) begin
          coeffs_294 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_295 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h127 == rs2[9:0]) begin
          coeffs_295 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_296 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h128 == rs2[9:0]) begin
          coeffs_296 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_297 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h129 == rs2[9:0]) begin
          coeffs_297 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_298 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h12a == rs2[9:0]) begin
          coeffs_298 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_299 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h12b == rs2[9:0]) begin
          coeffs_299 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_300 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h12c == rs2[9:0]) begin
          coeffs_300 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_301 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h12d == rs2[9:0]) begin
          coeffs_301 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_302 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h12e == rs2[9:0]) begin
          coeffs_302 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_303 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h12f == rs2[9:0]) begin
          coeffs_303 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_304 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h130 == rs2[9:0]) begin
          coeffs_304 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_305 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h131 == rs2[9:0]) begin
          coeffs_305 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_306 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h132 == rs2[9:0]) begin
          coeffs_306 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_307 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h133 == rs2[9:0]) begin
          coeffs_307 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_308 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h134 == rs2[9:0]) begin
          coeffs_308 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_309 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h135 == rs2[9:0]) begin
          coeffs_309 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_310 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h136 == rs2[9:0]) begin
          coeffs_310 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_311 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h137 == rs2[9:0]) begin
          coeffs_311 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_312 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h138 == rs2[9:0]) begin
          coeffs_312 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_313 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h139 == rs2[9:0]) begin
          coeffs_313 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_314 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h13a == rs2[9:0]) begin
          coeffs_314 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_315 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h13b == rs2[9:0]) begin
          coeffs_315 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_316 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h13c == rs2[9:0]) begin
          coeffs_316 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_317 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h13d == rs2[9:0]) begin
          coeffs_317 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_318 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h13e == rs2[9:0]) begin
          coeffs_318 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_319 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h13f == rs2[9:0]) begin
          coeffs_319 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_320 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h140 == rs2[9:0]) begin
          coeffs_320 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_321 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h141 == rs2[9:0]) begin
          coeffs_321 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_322 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h142 == rs2[9:0]) begin
          coeffs_322 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_323 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h143 == rs2[9:0]) begin
          coeffs_323 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_324 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h144 == rs2[9:0]) begin
          coeffs_324 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_325 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h145 == rs2[9:0]) begin
          coeffs_325 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_326 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h146 == rs2[9:0]) begin
          coeffs_326 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_327 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h147 == rs2[9:0]) begin
          coeffs_327 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_328 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h148 == rs2[9:0]) begin
          coeffs_328 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_329 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h149 == rs2[9:0]) begin
          coeffs_329 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_330 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h14a == rs2[9:0]) begin
          coeffs_330 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_331 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h14b == rs2[9:0]) begin
          coeffs_331 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_332 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h14c == rs2[9:0]) begin
          coeffs_332 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_333 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h14d == rs2[9:0]) begin
          coeffs_333 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_334 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h14e == rs2[9:0]) begin
          coeffs_334 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_335 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h14f == rs2[9:0]) begin
          coeffs_335 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_336 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h150 == rs2[9:0]) begin
          coeffs_336 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_337 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h151 == rs2[9:0]) begin
          coeffs_337 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_338 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h152 == rs2[9:0]) begin
          coeffs_338 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_339 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h153 == rs2[9:0]) begin
          coeffs_339 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_340 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h154 == rs2[9:0]) begin
          coeffs_340 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_341 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h155 == rs2[9:0]) begin
          coeffs_341 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_342 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h156 == rs2[9:0]) begin
          coeffs_342 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_343 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h157 == rs2[9:0]) begin
          coeffs_343 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_344 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h158 == rs2[9:0]) begin
          coeffs_344 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_345 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h159 == rs2[9:0]) begin
          coeffs_345 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_346 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h15a == rs2[9:0]) begin
          coeffs_346 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_347 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h15b == rs2[9:0]) begin
          coeffs_347 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_348 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h15c == rs2[9:0]) begin
          coeffs_348 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_349 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h15d == rs2[9:0]) begin
          coeffs_349 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_350 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h15e == rs2[9:0]) begin
          coeffs_350 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_351 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h15f == rs2[9:0]) begin
          coeffs_351 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_352 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h160 == rs2[9:0]) begin
          coeffs_352 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_353 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h161 == rs2[9:0]) begin
          coeffs_353 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_354 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h162 == rs2[9:0]) begin
          coeffs_354 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_355 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h163 == rs2[9:0]) begin
          coeffs_355 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_356 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h164 == rs2[9:0]) begin
          coeffs_356 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_357 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h165 == rs2[9:0]) begin
          coeffs_357 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_358 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h166 == rs2[9:0]) begin
          coeffs_358 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_359 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h167 == rs2[9:0]) begin
          coeffs_359 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_360 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h168 == rs2[9:0]) begin
          coeffs_360 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_361 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h169 == rs2[9:0]) begin
          coeffs_361 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_362 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h16a == rs2[9:0]) begin
          coeffs_362 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_363 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h16b == rs2[9:0]) begin
          coeffs_363 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_364 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h16c == rs2[9:0]) begin
          coeffs_364 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_365 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h16d == rs2[9:0]) begin
          coeffs_365 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_366 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h16e == rs2[9:0]) begin
          coeffs_366 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_367 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h16f == rs2[9:0]) begin
          coeffs_367 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_368 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h170 == rs2[9:0]) begin
          coeffs_368 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_369 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h171 == rs2[9:0]) begin
          coeffs_369 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_370 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h172 == rs2[9:0]) begin
          coeffs_370 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_371 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h173 == rs2[9:0]) begin
          coeffs_371 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_372 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h174 == rs2[9:0]) begin
          coeffs_372 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_373 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h175 == rs2[9:0]) begin
          coeffs_373 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_374 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h176 == rs2[9:0]) begin
          coeffs_374 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_375 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h177 == rs2[9:0]) begin
          coeffs_375 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_376 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h178 == rs2[9:0]) begin
          coeffs_376 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_377 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h179 == rs2[9:0]) begin
          coeffs_377 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_378 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h17a == rs2[9:0]) begin
          coeffs_378 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_379 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h17b == rs2[9:0]) begin
          coeffs_379 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_380 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h17c == rs2[9:0]) begin
          coeffs_380 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_381 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h17d == rs2[9:0]) begin
          coeffs_381 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_382 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h17e == rs2[9:0]) begin
          coeffs_382 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_383 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h17f == rs2[9:0]) begin
          coeffs_383 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_384 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h180 == rs2[9:0]) begin
          coeffs_384 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_385 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h181 == rs2[9:0]) begin
          coeffs_385 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_386 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h182 == rs2[9:0]) begin
          coeffs_386 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_387 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h183 == rs2[9:0]) begin
          coeffs_387 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_388 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h184 == rs2[9:0]) begin
          coeffs_388 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_389 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h185 == rs2[9:0]) begin
          coeffs_389 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_390 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h186 == rs2[9:0]) begin
          coeffs_390 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_391 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h187 == rs2[9:0]) begin
          coeffs_391 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_392 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h188 == rs2[9:0]) begin
          coeffs_392 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_393 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h189 == rs2[9:0]) begin
          coeffs_393 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_394 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h18a == rs2[9:0]) begin
          coeffs_394 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_395 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h18b == rs2[9:0]) begin
          coeffs_395 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_396 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h18c == rs2[9:0]) begin
          coeffs_396 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_397 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h18d == rs2[9:0]) begin
          coeffs_397 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_398 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h18e == rs2[9:0]) begin
          coeffs_398 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_399 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h18f == rs2[9:0]) begin
          coeffs_399 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_400 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h190 == rs2[9:0]) begin
          coeffs_400 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_401 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h191 == rs2[9:0]) begin
          coeffs_401 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_402 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h192 == rs2[9:0]) begin
          coeffs_402 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_403 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h193 == rs2[9:0]) begin
          coeffs_403 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_404 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h194 == rs2[9:0]) begin
          coeffs_404 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_405 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h195 == rs2[9:0]) begin
          coeffs_405 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_406 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h196 == rs2[9:0]) begin
          coeffs_406 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_407 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h197 == rs2[9:0]) begin
          coeffs_407 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_408 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h198 == rs2[9:0]) begin
          coeffs_408 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_409 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h199 == rs2[9:0]) begin
          coeffs_409 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_410 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h19a == rs2[9:0]) begin
          coeffs_410 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_411 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h19b == rs2[9:0]) begin
          coeffs_411 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_412 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h19c == rs2[9:0]) begin
          coeffs_412 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_413 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h19d == rs2[9:0]) begin
          coeffs_413 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_414 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h19e == rs2[9:0]) begin
          coeffs_414 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_415 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h19f == rs2[9:0]) begin
          coeffs_415 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_416 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a0 == rs2[9:0]) begin
          coeffs_416 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_417 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a1 == rs2[9:0]) begin
          coeffs_417 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_418 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a2 == rs2[9:0]) begin
          coeffs_418 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_419 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a3 == rs2[9:0]) begin
          coeffs_419 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_420 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a4 == rs2[9:0]) begin
          coeffs_420 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_421 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a5 == rs2[9:0]) begin
          coeffs_421 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_422 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a6 == rs2[9:0]) begin
          coeffs_422 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_423 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a7 == rs2[9:0]) begin
          coeffs_423 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_424 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a8 == rs2[9:0]) begin
          coeffs_424 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_425 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a9 == rs2[9:0]) begin
          coeffs_425 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_426 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1aa == rs2[9:0]) begin
          coeffs_426 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_427 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ab == rs2[9:0]) begin
          coeffs_427 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_428 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ac == rs2[9:0]) begin
          coeffs_428 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_429 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ad == rs2[9:0]) begin
          coeffs_429 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_430 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ae == rs2[9:0]) begin
          coeffs_430 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_431 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1af == rs2[9:0]) begin
          coeffs_431 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_432 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b0 == rs2[9:0]) begin
          coeffs_432 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_433 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b1 == rs2[9:0]) begin
          coeffs_433 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_434 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b2 == rs2[9:0]) begin
          coeffs_434 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_435 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b3 == rs2[9:0]) begin
          coeffs_435 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_436 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b4 == rs2[9:0]) begin
          coeffs_436 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_437 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b5 == rs2[9:0]) begin
          coeffs_437 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_438 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b6 == rs2[9:0]) begin
          coeffs_438 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_439 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b7 == rs2[9:0]) begin
          coeffs_439 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_440 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b8 == rs2[9:0]) begin
          coeffs_440 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_441 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b9 == rs2[9:0]) begin
          coeffs_441 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_442 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ba == rs2[9:0]) begin
          coeffs_442 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_443 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1bb == rs2[9:0]) begin
          coeffs_443 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_444 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1bc == rs2[9:0]) begin
          coeffs_444 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_445 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1bd == rs2[9:0]) begin
          coeffs_445 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_446 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1be == rs2[9:0]) begin
          coeffs_446 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_447 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1bf == rs2[9:0]) begin
          coeffs_447 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_448 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c0 == rs2[9:0]) begin
          coeffs_448 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_449 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c1 == rs2[9:0]) begin
          coeffs_449 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_450 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c2 == rs2[9:0]) begin
          coeffs_450 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_451 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c3 == rs2[9:0]) begin
          coeffs_451 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_452 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c4 == rs2[9:0]) begin
          coeffs_452 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_453 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c5 == rs2[9:0]) begin
          coeffs_453 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_454 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c6 == rs2[9:0]) begin
          coeffs_454 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_455 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c7 == rs2[9:0]) begin
          coeffs_455 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_456 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c8 == rs2[9:0]) begin
          coeffs_456 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_457 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c9 == rs2[9:0]) begin
          coeffs_457 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_458 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ca == rs2[9:0]) begin
          coeffs_458 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_459 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1cb == rs2[9:0]) begin
          coeffs_459 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_460 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1cc == rs2[9:0]) begin
          coeffs_460 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_461 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1cd == rs2[9:0]) begin
          coeffs_461 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_462 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ce == rs2[9:0]) begin
          coeffs_462 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_463 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1cf == rs2[9:0]) begin
          coeffs_463 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_464 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d0 == rs2[9:0]) begin
          coeffs_464 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_465 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d1 == rs2[9:0]) begin
          coeffs_465 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_466 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d2 == rs2[9:0]) begin
          coeffs_466 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_467 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d3 == rs2[9:0]) begin
          coeffs_467 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_468 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d4 == rs2[9:0]) begin
          coeffs_468 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_469 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d5 == rs2[9:0]) begin
          coeffs_469 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_470 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d6 == rs2[9:0]) begin
          coeffs_470 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_471 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d7 == rs2[9:0]) begin
          coeffs_471 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_472 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d8 == rs2[9:0]) begin
          coeffs_472 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_473 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d9 == rs2[9:0]) begin
          coeffs_473 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_474 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1da == rs2[9:0]) begin
          coeffs_474 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_475 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1db == rs2[9:0]) begin
          coeffs_475 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_476 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1dc == rs2[9:0]) begin
          coeffs_476 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_477 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1dd == rs2[9:0]) begin
          coeffs_477 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_478 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1de == rs2[9:0]) begin
          coeffs_478 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_479 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1df == rs2[9:0]) begin
          coeffs_479 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_480 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e0 == rs2[9:0]) begin
          coeffs_480 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_481 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e1 == rs2[9:0]) begin
          coeffs_481 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_482 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e2 == rs2[9:0]) begin
          coeffs_482 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_483 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e3 == rs2[9:0]) begin
          coeffs_483 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_484 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e4 == rs2[9:0]) begin
          coeffs_484 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_485 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e5 == rs2[9:0]) begin
          coeffs_485 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_486 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e6 == rs2[9:0]) begin
          coeffs_486 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_487 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e7 == rs2[9:0]) begin
          coeffs_487 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_488 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e8 == rs2[9:0]) begin
          coeffs_488 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_489 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e9 == rs2[9:0]) begin
          coeffs_489 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_490 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ea == rs2[9:0]) begin
          coeffs_490 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_491 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1eb == rs2[9:0]) begin
          coeffs_491 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_492 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ec == rs2[9:0]) begin
          coeffs_492 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_493 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ed == rs2[9:0]) begin
          coeffs_493 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_494 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ee == rs2[9:0]) begin
          coeffs_494 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_495 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ef == rs2[9:0]) begin
          coeffs_495 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_496 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f0 == rs2[9:0]) begin
          coeffs_496 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_497 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f1 == rs2[9:0]) begin
          coeffs_497 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_498 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f2 == rs2[9:0]) begin
          coeffs_498 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_499 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f3 == rs2[9:0]) begin
          coeffs_499 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_500 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f4 == rs2[9:0]) begin
          coeffs_500 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_501 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f5 == rs2[9:0]) begin
          coeffs_501 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_502 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f6 == rs2[9:0]) begin
          coeffs_502 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_503 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f7 == rs2[9:0]) begin
          coeffs_503 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_504 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f8 == rs2[9:0]) begin
          coeffs_504 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_505 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f9 == rs2[9:0]) begin
          coeffs_505 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_506 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1fa == rs2[9:0]) begin
          coeffs_506 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_507 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1fb == rs2[9:0]) begin
          coeffs_507 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_508 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1fc == rs2[9:0]) begin
          coeffs_508 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_509 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1fd == rs2[9:0]) begin
          coeffs_509 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_510 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1fe == rs2[9:0]) begin
          coeffs_510 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_511 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ff == rs2[9:0]) begin
          coeffs_511 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_512 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h200 == rs2[9:0]) begin
          coeffs_512 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_513 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h201 == rs2[9:0]) begin
          coeffs_513 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_514 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h202 == rs2[9:0]) begin
          coeffs_514 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_515 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h203 == rs2[9:0]) begin
          coeffs_515 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_516 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h204 == rs2[9:0]) begin
          coeffs_516 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_517 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h205 == rs2[9:0]) begin
          coeffs_517 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_518 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h206 == rs2[9:0]) begin
          coeffs_518 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_519 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h207 == rs2[9:0]) begin
          coeffs_519 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_520 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h208 == rs2[9:0]) begin
          coeffs_520 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_521 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h209 == rs2[9:0]) begin
          coeffs_521 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_522 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h20a == rs2[9:0]) begin
          coeffs_522 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_523 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h20b == rs2[9:0]) begin
          coeffs_523 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_524 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h20c == rs2[9:0]) begin
          coeffs_524 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_525 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h20d == rs2[9:0]) begin
          coeffs_525 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_526 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h20e == rs2[9:0]) begin
          coeffs_526 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_527 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h20f == rs2[9:0]) begin
          coeffs_527 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_528 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h210 == rs2[9:0]) begin
          coeffs_528 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_529 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h211 == rs2[9:0]) begin
          coeffs_529 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_530 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h212 == rs2[9:0]) begin
          coeffs_530 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_531 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h213 == rs2[9:0]) begin
          coeffs_531 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_532 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h214 == rs2[9:0]) begin
          coeffs_532 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_533 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h215 == rs2[9:0]) begin
          coeffs_533 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_534 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h216 == rs2[9:0]) begin
          coeffs_534 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_535 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h217 == rs2[9:0]) begin
          coeffs_535 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_536 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h218 == rs2[9:0]) begin
          coeffs_536 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_537 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h219 == rs2[9:0]) begin
          coeffs_537 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_538 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h21a == rs2[9:0]) begin
          coeffs_538 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_539 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h21b == rs2[9:0]) begin
          coeffs_539 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_540 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h21c == rs2[9:0]) begin
          coeffs_540 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_541 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h21d == rs2[9:0]) begin
          coeffs_541 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_542 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h21e == rs2[9:0]) begin
          coeffs_542 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_543 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h21f == rs2[9:0]) begin
          coeffs_543 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_544 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h220 == rs2[9:0]) begin
          coeffs_544 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_545 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h221 == rs2[9:0]) begin
          coeffs_545 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_546 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h222 == rs2[9:0]) begin
          coeffs_546 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_547 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h223 == rs2[9:0]) begin
          coeffs_547 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_548 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h224 == rs2[9:0]) begin
          coeffs_548 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_549 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h225 == rs2[9:0]) begin
          coeffs_549 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_550 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h226 == rs2[9:0]) begin
          coeffs_550 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_551 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h227 == rs2[9:0]) begin
          coeffs_551 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_552 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h228 == rs2[9:0]) begin
          coeffs_552 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_553 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h229 == rs2[9:0]) begin
          coeffs_553 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_554 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h22a == rs2[9:0]) begin
          coeffs_554 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_555 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h22b == rs2[9:0]) begin
          coeffs_555 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_556 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h22c == rs2[9:0]) begin
          coeffs_556 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_557 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h22d == rs2[9:0]) begin
          coeffs_557 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_558 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h22e == rs2[9:0]) begin
          coeffs_558 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_559 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h22f == rs2[9:0]) begin
          coeffs_559 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_560 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h230 == rs2[9:0]) begin
          coeffs_560 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_561 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h231 == rs2[9:0]) begin
          coeffs_561 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_562 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h232 == rs2[9:0]) begin
          coeffs_562 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_563 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h233 == rs2[9:0]) begin
          coeffs_563 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_564 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h234 == rs2[9:0]) begin
          coeffs_564 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_565 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h235 == rs2[9:0]) begin
          coeffs_565 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_566 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h236 == rs2[9:0]) begin
          coeffs_566 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_567 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h237 == rs2[9:0]) begin
          coeffs_567 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_568 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h238 == rs2[9:0]) begin
          coeffs_568 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_569 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h239 == rs2[9:0]) begin
          coeffs_569 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_570 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h23a == rs2[9:0]) begin
          coeffs_570 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_571 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h23b == rs2[9:0]) begin
          coeffs_571 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_572 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h23c == rs2[9:0]) begin
          coeffs_572 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_573 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h23d == rs2[9:0]) begin
          coeffs_573 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_574 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h23e == rs2[9:0]) begin
          coeffs_574 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_575 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h23f == rs2[9:0]) begin
          coeffs_575 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_576 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h240 == rs2[9:0]) begin
          coeffs_576 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_577 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h241 == rs2[9:0]) begin
          coeffs_577 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_578 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h242 == rs2[9:0]) begin
          coeffs_578 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_579 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h243 == rs2[9:0]) begin
          coeffs_579 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_580 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h244 == rs2[9:0]) begin
          coeffs_580 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_581 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h245 == rs2[9:0]) begin
          coeffs_581 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_582 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h246 == rs2[9:0]) begin
          coeffs_582 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_583 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h247 == rs2[9:0]) begin
          coeffs_583 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_584 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h248 == rs2[9:0]) begin
          coeffs_584 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_585 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h249 == rs2[9:0]) begin
          coeffs_585 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_586 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h24a == rs2[9:0]) begin
          coeffs_586 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_587 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h24b == rs2[9:0]) begin
          coeffs_587 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_588 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h24c == rs2[9:0]) begin
          coeffs_588 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_589 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h24d == rs2[9:0]) begin
          coeffs_589 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_590 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h24e == rs2[9:0]) begin
          coeffs_590 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_591 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h24f == rs2[9:0]) begin
          coeffs_591 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_592 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h250 == rs2[9:0]) begin
          coeffs_592 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_593 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h251 == rs2[9:0]) begin
          coeffs_593 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_594 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h252 == rs2[9:0]) begin
          coeffs_594 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_595 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h253 == rs2[9:0]) begin
          coeffs_595 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_596 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h254 == rs2[9:0]) begin
          coeffs_596 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_597 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h255 == rs2[9:0]) begin
          coeffs_597 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_598 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h256 == rs2[9:0]) begin
          coeffs_598 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_599 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h257 == rs2[9:0]) begin
          coeffs_599 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_600 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h258 == rs2[9:0]) begin
          coeffs_600 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_601 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h259 == rs2[9:0]) begin
          coeffs_601 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_602 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h25a == rs2[9:0]) begin
          coeffs_602 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_603 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h25b == rs2[9:0]) begin
          coeffs_603 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_604 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h25c == rs2[9:0]) begin
          coeffs_604 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_605 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h25d == rs2[9:0]) begin
          coeffs_605 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_606 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h25e == rs2[9:0]) begin
          coeffs_606 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_607 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h25f == rs2[9:0]) begin
          coeffs_607 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_608 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h260 == rs2[9:0]) begin
          coeffs_608 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_609 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h261 == rs2[9:0]) begin
          coeffs_609 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_610 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h262 == rs2[9:0]) begin
          coeffs_610 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_611 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h263 == rs2[9:0]) begin
          coeffs_611 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_612 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h264 == rs2[9:0]) begin
          coeffs_612 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_613 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h265 == rs2[9:0]) begin
          coeffs_613 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_614 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h266 == rs2[9:0]) begin
          coeffs_614 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_615 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h267 == rs2[9:0]) begin
          coeffs_615 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_616 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h268 == rs2[9:0]) begin
          coeffs_616 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_617 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h269 == rs2[9:0]) begin
          coeffs_617 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_618 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h26a == rs2[9:0]) begin
          coeffs_618 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_619 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h26b == rs2[9:0]) begin
          coeffs_619 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_620 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h26c == rs2[9:0]) begin
          coeffs_620 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_621 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h26d == rs2[9:0]) begin
          coeffs_621 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_622 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h26e == rs2[9:0]) begin
          coeffs_622 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_623 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h26f == rs2[9:0]) begin
          coeffs_623 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_624 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h270 == rs2[9:0]) begin
          coeffs_624 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_625 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h271 == rs2[9:0]) begin
          coeffs_625 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_626 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h272 == rs2[9:0]) begin
          coeffs_626 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_627 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h273 == rs2[9:0]) begin
          coeffs_627 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_628 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h274 == rs2[9:0]) begin
          coeffs_628 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_629 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h275 == rs2[9:0]) begin
          coeffs_629 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_630 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h276 == rs2[9:0]) begin
          coeffs_630 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_631 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h277 == rs2[9:0]) begin
          coeffs_631 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_632 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h278 == rs2[9:0]) begin
          coeffs_632 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_633 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h279 == rs2[9:0]) begin
          coeffs_633 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_634 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h27a == rs2[9:0]) begin
          coeffs_634 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_635 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h27b == rs2[9:0]) begin
          coeffs_635 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_636 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h27c == rs2[9:0]) begin
          coeffs_636 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_637 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h27d == rs2[9:0]) begin
          coeffs_637 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_638 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h27e == rs2[9:0]) begin
          coeffs_638 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_639 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h27f == rs2[9:0]) begin
          coeffs_639 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_640 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h280 == rs2[9:0]) begin
          coeffs_640 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_641 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h281 == rs2[9:0]) begin
          coeffs_641 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_642 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h282 == rs2[9:0]) begin
          coeffs_642 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_643 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h283 == rs2[9:0]) begin
          coeffs_643 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_644 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h284 == rs2[9:0]) begin
          coeffs_644 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_645 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h285 == rs2[9:0]) begin
          coeffs_645 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_646 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h286 == rs2[9:0]) begin
          coeffs_646 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_647 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h287 == rs2[9:0]) begin
          coeffs_647 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_648 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h288 == rs2[9:0]) begin
          coeffs_648 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_649 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h289 == rs2[9:0]) begin
          coeffs_649 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_650 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h28a == rs2[9:0]) begin
          coeffs_650 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_651 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h28b == rs2[9:0]) begin
          coeffs_651 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_652 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h28c == rs2[9:0]) begin
          coeffs_652 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_653 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h28d == rs2[9:0]) begin
          coeffs_653 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_654 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h28e == rs2[9:0]) begin
          coeffs_654 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_655 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h28f == rs2[9:0]) begin
          coeffs_655 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_656 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h290 == rs2[9:0]) begin
          coeffs_656 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_657 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h291 == rs2[9:0]) begin
          coeffs_657 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_658 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h292 == rs2[9:0]) begin
          coeffs_658 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_659 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h293 == rs2[9:0]) begin
          coeffs_659 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_660 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h294 == rs2[9:0]) begin
          coeffs_660 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_661 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h295 == rs2[9:0]) begin
          coeffs_661 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_662 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h296 == rs2[9:0]) begin
          coeffs_662 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_663 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h297 == rs2[9:0]) begin
          coeffs_663 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_664 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h298 == rs2[9:0]) begin
          coeffs_664 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_665 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h299 == rs2[9:0]) begin
          coeffs_665 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_666 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h29a == rs2[9:0]) begin
          coeffs_666 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_667 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h29b == rs2[9:0]) begin
          coeffs_667 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_668 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h29c == rs2[9:0]) begin
          coeffs_668 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_669 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h29d == rs2[9:0]) begin
          coeffs_669 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_670 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h29e == rs2[9:0]) begin
          coeffs_670 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_671 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h29f == rs2[9:0]) begin
          coeffs_671 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_672 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a0 == rs2[9:0]) begin
          coeffs_672 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_673 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a1 == rs2[9:0]) begin
          coeffs_673 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_674 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a2 == rs2[9:0]) begin
          coeffs_674 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_675 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a3 == rs2[9:0]) begin
          coeffs_675 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_676 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a4 == rs2[9:0]) begin
          coeffs_676 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_677 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a5 == rs2[9:0]) begin
          coeffs_677 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_678 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a6 == rs2[9:0]) begin
          coeffs_678 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_679 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a7 == rs2[9:0]) begin
          coeffs_679 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_680 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a8 == rs2[9:0]) begin
          coeffs_680 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_681 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a9 == rs2[9:0]) begin
          coeffs_681 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_682 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2aa == rs2[9:0]) begin
          coeffs_682 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_683 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ab == rs2[9:0]) begin
          coeffs_683 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_684 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ac == rs2[9:0]) begin
          coeffs_684 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_685 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ad == rs2[9:0]) begin
          coeffs_685 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_686 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ae == rs2[9:0]) begin
          coeffs_686 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_687 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2af == rs2[9:0]) begin
          coeffs_687 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_688 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b0 == rs2[9:0]) begin
          coeffs_688 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_689 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b1 == rs2[9:0]) begin
          coeffs_689 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_690 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b2 == rs2[9:0]) begin
          coeffs_690 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_691 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b3 == rs2[9:0]) begin
          coeffs_691 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_692 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b4 == rs2[9:0]) begin
          coeffs_692 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_693 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b5 == rs2[9:0]) begin
          coeffs_693 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_694 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b6 == rs2[9:0]) begin
          coeffs_694 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_695 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b7 == rs2[9:0]) begin
          coeffs_695 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_696 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b8 == rs2[9:0]) begin
          coeffs_696 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_697 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b9 == rs2[9:0]) begin
          coeffs_697 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_698 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ba == rs2[9:0]) begin
          coeffs_698 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_699 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2bb == rs2[9:0]) begin
          coeffs_699 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_700 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2bc == rs2[9:0]) begin
          coeffs_700 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_701 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2bd == rs2[9:0]) begin
          coeffs_701 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_702 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2be == rs2[9:0]) begin
          coeffs_702 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_703 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2bf == rs2[9:0]) begin
          coeffs_703 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_704 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c0 == rs2[9:0]) begin
          coeffs_704 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_705 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c1 == rs2[9:0]) begin
          coeffs_705 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_706 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c2 == rs2[9:0]) begin
          coeffs_706 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_707 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c3 == rs2[9:0]) begin
          coeffs_707 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_708 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c4 == rs2[9:0]) begin
          coeffs_708 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_709 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c5 == rs2[9:0]) begin
          coeffs_709 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_710 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c6 == rs2[9:0]) begin
          coeffs_710 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_711 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c7 == rs2[9:0]) begin
          coeffs_711 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_712 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c8 == rs2[9:0]) begin
          coeffs_712 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_713 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c9 == rs2[9:0]) begin
          coeffs_713 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_714 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ca == rs2[9:0]) begin
          coeffs_714 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_715 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2cb == rs2[9:0]) begin
          coeffs_715 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_716 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2cc == rs2[9:0]) begin
          coeffs_716 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_717 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2cd == rs2[9:0]) begin
          coeffs_717 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_718 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ce == rs2[9:0]) begin
          coeffs_718 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_719 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2cf == rs2[9:0]) begin
          coeffs_719 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_720 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d0 == rs2[9:0]) begin
          coeffs_720 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_721 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d1 == rs2[9:0]) begin
          coeffs_721 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_722 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d2 == rs2[9:0]) begin
          coeffs_722 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_723 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d3 == rs2[9:0]) begin
          coeffs_723 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_724 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d4 == rs2[9:0]) begin
          coeffs_724 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_725 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d5 == rs2[9:0]) begin
          coeffs_725 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_726 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d6 == rs2[9:0]) begin
          coeffs_726 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_727 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d7 == rs2[9:0]) begin
          coeffs_727 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_728 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d8 == rs2[9:0]) begin
          coeffs_728 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_729 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d9 == rs2[9:0]) begin
          coeffs_729 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_730 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2da == rs2[9:0]) begin
          coeffs_730 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_731 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2db == rs2[9:0]) begin
          coeffs_731 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_732 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2dc == rs2[9:0]) begin
          coeffs_732 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_733 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2dd == rs2[9:0]) begin
          coeffs_733 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_734 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2de == rs2[9:0]) begin
          coeffs_734 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_735 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2df == rs2[9:0]) begin
          coeffs_735 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_736 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e0 == rs2[9:0]) begin
          coeffs_736 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_737 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e1 == rs2[9:0]) begin
          coeffs_737 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_738 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e2 == rs2[9:0]) begin
          coeffs_738 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_739 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e3 == rs2[9:0]) begin
          coeffs_739 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_740 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e4 == rs2[9:0]) begin
          coeffs_740 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_741 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e5 == rs2[9:0]) begin
          coeffs_741 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_742 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e6 == rs2[9:0]) begin
          coeffs_742 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_743 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e7 == rs2[9:0]) begin
          coeffs_743 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_744 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e8 == rs2[9:0]) begin
          coeffs_744 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_745 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e9 == rs2[9:0]) begin
          coeffs_745 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_746 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ea == rs2[9:0]) begin
          coeffs_746 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_747 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2eb == rs2[9:0]) begin
          coeffs_747 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_748 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ec == rs2[9:0]) begin
          coeffs_748 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_749 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ed == rs2[9:0]) begin
          coeffs_749 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_750 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ee == rs2[9:0]) begin
          coeffs_750 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_751 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ef == rs2[9:0]) begin
          coeffs_751 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_752 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f0 == rs2[9:0]) begin
          coeffs_752 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_753 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f1 == rs2[9:0]) begin
          coeffs_753 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_754 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f2 == rs2[9:0]) begin
          coeffs_754 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_755 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f3 == rs2[9:0]) begin
          coeffs_755 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_756 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f4 == rs2[9:0]) begin
          coeffs_756 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_757 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f5 == rs2[9:0]) begin
          coeffs_757 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_758 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f6 == rs2[9:0]) begin
          coeffs_758 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_759 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f7 == rs2[9:0]) begin
          coeffs_759 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_760 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f8 == rs2[9:0]) begin
          coeffs_760 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_761 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f9 == rs2[9:0]) begin
          coeffs_761 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_762 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2fa == rs2[9:0]) begin
          coeffs_762 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_763 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2fb == rs2[9:0]) begin
          coeffs_763 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_764 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2fc == rs2[9:0]) begin
          coeffs_764 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_765 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2fd == rs2[9:0]) begin
          coeffs_765 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_766 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2fe == rs2[9:0]) begin
          coeffs_766 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_767 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ff == rs2[9:0]) begin
          coeffs_767 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_768 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h300 == rs2[9:0]) begin
          coeffs_768 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_769 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h301 == rs2[9:0]) begin
          coeffs_769 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_770 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h302 == rs2[9:0]) begin
          coeffs_770 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_771 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h303 == rs2[9:0]) begin
          coeffs_771 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_772 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h304 == rs2[9:0]) begin
          coeffs_772 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_773 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h305 == rs2[9:0]) begin
          coeffs_773 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_774 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h306 == rs2[9:0]) begin
          coeffs_774 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_775 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h307 == rs2[9:0]) begin
          coeffs_775 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_776 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h308 == rs2[9:0]) begin
          coeffs_776 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_777 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h309 == rs2[9:0]) begin
          coeffs_777 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_778 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h30a == rs2[9:0]) begin
          coeffs_778 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_779 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h30b == rs2[9:0]) begin
          coeffs_779 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_780 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h30c == rs2[9:0]) begin
          coeffs_780 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_781 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h30d == rs2[9:0]) begin
          coeffs_781 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_782 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h30e == rs2[9:0]) begin
          coeffs_782 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_783 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h30f == rs2[9:0]) begin
          coeffs_783 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_784 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h310 == rs2[9:0]) begin
          coeffs_784 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_785 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h311 == rs2[9:0]) begin
          coeffs_785 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_786 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h312 == rs2[9:0]) begin
          coeffs_786 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_787 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h313 == rs2[9:0]) begin
          coeffs_787 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_788 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h314 == rs2[9:0]) begin
          coeffs_788 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_789 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h315 == rs2[9:0]) begin
          coeffs_789 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_790 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h316 == rs2[9:0]) begin
          coeffs_790 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_791 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h317 == rs2[9:0]) begin
          coeffs_791 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_792 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h318 == rs2[9:0]) begin
          coeffs_792 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_793 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h319 == rs2[9:0]) begin
          coeffs_793 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_794 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h31a == rs2[9:0]) begin
          coeffs_794 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_795 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h31b == rs2[9:0]) begin
          coeffs_795 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_796 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h31c == rs2[9:0]) begin
          coeffs_796 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_797 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h31d == rs2[9:0]) begin
          coeffs_797 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_798 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h31e == rs2[9:0]) begin
          coeffs_798 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_799 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h31f == rs2[9:0]) begin
          coeffs_799 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_800 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h320 == rs2[9:0]) begin
          coeffs_800 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_801 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h321 == rs2[9:0]) begin
          coeffs_801 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_802 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h322 == rs2[9:0]) begin
          coeffs_802 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_803 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h323 == rs2[9:0]) begin
          coeffs_803 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_804 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h324 == rs2[9:0]) begin
          coeffs_804 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_805 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h325 == rs2[9:0]) begin
          coeffs_805 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_806 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h326 == rs2[9:0]) begin
          coeffs_806 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_807 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h327 == rs2[9:0]) begin
          coeffs_807 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_808 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h328 == rs2[9:0]) begin
          coeffs_808 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_809 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h329 == rs2[9:0]) begin
          coeffs_809 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_810 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h32a == rs2[9:0]) begin
          coeffs_810 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_811 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h32b == rs2[9:0]) begin
          coeffs_811 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_812 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h32c == rs2[9:0]) begin
          coeffs_812 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_813 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h32d == rs2[9:0]) begin
          coeffs_813 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_814 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h32e == rs2[9:0]) begin
          coeffs_814 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_815 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h32f == rs2[9:0]) begin
          coeffs_815 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_816 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h330 == rs2[9:0]) begin
          coeffs_816 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_817 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h331 == rs2[9:0]) begin
          coeffs_817 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_818 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h332 == rs2[9:0]) begin
          coeffs_818 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_819 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h333 == rs2[9:0]) begin
          coeffs_819 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_820 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h334 == rs2[9:0]) begin
          coeffs_820 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_821 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h335 == rs2[9:0]) begin
          coeffs_821 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_822 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h336 == rs2[9:0]) begin
          coeffs_822 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_823 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h337 == rs2[9:0]) begin
          coeffs_823 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_824 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h338 == rs2[9:0]) begin
          coeffs_824 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_825 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h339 == rs2[9:0]) begin
          coeffs_825 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_826 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h33a == rs2[9:0]) begin
          coeffs_826 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_827 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h33b == rs2[9:0]) begin
          coeffs_827 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_828 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h33c == rs2[9:0]) begin
          coeffs_828 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_829 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h33d == rs2[9:0]) begin
          coeffs_829 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_830 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h33e == rs2[9:0]) begin
          coeffs_830 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_831 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h33f == rs2[9:0]) begin
          coeffs_831 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_832 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h340 == rs2[9:0]) begin
          coeffs_832 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_833 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h341 == rs2[9:0]) begin
          coeffs_833 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_834 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h342 == rs2[9:0]) begin
          coeffs_834 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_835 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h343 == rs2[9:0]) begin
          coeffs_835 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_836 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h344 == rs2[9:0]) begin
          coeffs_836 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_837 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h345 == rs2[9:0]) begin
          coeffs_837 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_838 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h346 == rs2[9:0]) begin
          coeffs_838 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_839 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h347 == rs2[9:0]) begin
          coeffs_839 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_840 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h348 == rs2[9:0]) begin
          coeffs_840 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_841 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h349 == rs2[9:0]) begin
          coeffs_841 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_842 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h34a == rs2[9:0]) begin
          coeffs_842 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_843 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h34b == rs2[9:0]) begin
          coeffs_843 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_844 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h34c == rs2[9:0]) begin
          coeffs_844 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_845 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h34d == rs2[9:0]) begin
          coeffs_845 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_846 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h34e == rs2[9:0]) begin
          coeffs_846 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_847 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h34f == rs2[9:0]) begin
          coeffs_847 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_848 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h350 == rs2[9:0]) begin
          coeffs_848 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_849 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h351 == rs2[9:0]) begin
          coeffs_849 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_850 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h352 == rs2[9:0]) begin
          coeffs_850 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_851 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h353 == rs2[9:0]) begin
          coeffs_851 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_852 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h354 == rs2[9:0]) begin
          coeffs_852 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_853 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h355 == rs2[9:0]) begin
          coeffs_853 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_854 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h356 == rs2[9:0]) begin
          coeffs_854 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_855 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h357 == rs2[9:0]) begin
          coeffs_855 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_856 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h358 == rs2[9:0]) begin
          coeffs_856 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_857 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h359 == rs2[9:0]) begin
          coeffs_857 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_858 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h35a == rs2[9:0]) begin
          coeffs_858 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_859 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h35b == rs2[9:0]) begin
          coeffs_859 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_860 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h35c == rs2[9:0]) begin
          coeffs_860 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_861 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h35d == rs2[9:0]) begin
          coeffs_861 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_862 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h35e == rs2[9:0]) begin
          coeffs_862 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_863 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h35f == rs2[9:0]) begin
          coeffs_863 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_864 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h360 == rs2[9:0]) begin
          coeffs_864 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_865 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h361 == rs2[9:0]) begin
          coeffs_865 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_866 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h362 == rs2[9:0]) begin
          coeffs_866 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_867 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h363 == rs2[9:0]) begin
          coeffs_867 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_868 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h364 == rs2[9:0]) begin
          coeffs_868 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_869 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h365 == rs2[9:0]) begin
          coeffs_869 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_870 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h366 == rs2[9:0]) begin
          coeffs_870 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_871 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h367 == rs2[9:0]) begin
          coeffs_871 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_872 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h368 == rs2[9:0]) begin
          coeffs_872 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_873 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h369 == rs2[9:0]) begin
          coeffs_873 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_874 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h36a == rs2[9:0]) begin
          coeffs_874 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_875 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h36b == rs2[9:0]) begin
          coeffs_875 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_876 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h36c == rs2[9:0]) begin
          coeffs_876 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_877 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h36d == rs2[9:0]) begin
          coeffs_877 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_878 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h36e == rs2[9:0]) begin
          coeffs_878 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_879 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h36f == rs2[9:0]) begin
          coeffs_879 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_880 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h370 == rs2[9:0]) begin
          coeffs_880 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_881 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h371 == rs2[9:0]) begin
          coeffs_881 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_882 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h372 == rs2[9:0]) begin
          coeffs_882 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_883 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h373 == rs2[9:0]) begin
          coeffs_883 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_884 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h374 == rs2[9:0]) begin
          coeffs_884 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_885 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h375 == rs2[9:0]) begin
          coeffs_885 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_886 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h376 == rs2[9:0]) begin
          coeffs_886 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_887 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h377 == rs2[9:0]) begin
          coeffs_887 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_888 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h378 == rs2[9:0]) begin
          coeffs_888 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_889 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h379 == rs2[9:0]) begin
          coeffs_889 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_890 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h37a == rs2[9:0]) begin
          coeffs_890 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_891 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h37b == rs2[9:0]) begin
          coeffs_891 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_892 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h37c == rs2[9:0]) begin
          coeffs_892 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_893 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h37d == rs2[9:0]) begin
          coeffs_893 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_894 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h37e == rs2[9:0]) begin
          coeffs_894 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_895 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h37f == rs2[9:0]) begin
          coeffs_895 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_896 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h380 == rs2[9:0]) begin
          coeffs_896 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_897 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h381 == rs2[9:0]) begin
          coeffs_897 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_898 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h382 == rs2[9:0]) begin
          coeffs_898 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_899 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h383 == rs2[9:0]) begin
          coeffs_899 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_900 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h384 == rs2[9:0]) begin
          coeffs_900 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_901 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h385 == rs2[9:0]) begin
          coeffs_901 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_902 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h386 == rs2[9:0]) begin
          coeffs_902 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_903 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h387 == rs2[9:0]) begin
          coeffs_903 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_904 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h388 == rs2[9:0]) begin
          coeffs_904 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_905 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h389 == rs2[9:0]) begin
          coeffs_905 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_906 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h38a == rs2[9:0]) begin
          coeffs_906 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_907 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h38b == rs2[9:0]) begin
          coeffs_907 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_908 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h38c == rs2[9:0]) begin
          coeffs_908 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_909 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h38d == rs2[9:0]) begin
          coeffs_909 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_910 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h38e == rs2[9:0]) begin
          coeffs_910 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_911 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h38f == rs2[9:0]) begin
          coeffs_911 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_912 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h390 == rs2[9:0]) begin
          coeffs_912 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_913 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h391 == rs2[9:0]) begin
          coeffs_913 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_914 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h392 == rs2[9:0]) begin
          coeffs_914 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_915 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h393 == rs2[9:0]) begin
          coeffs_915 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_916 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h394 == rs2[9:0]) begin
          coeffs_916 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_917 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h395 == rs2[9:0]) begin
          coeffs_917 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_918 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h396 == rs2[9:0]) begin
          coeffs_918 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_919 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h397 == rs2[9:0]) begin
          coeffs_919 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_920 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h398 == rs2[9:0]) begin
          coeffs_920 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_921 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h399 == rs2[9:0]) begin
          coeffs_921 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_922 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h39a == rs2[9:0]) begin
          coeffs_922 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_923 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h39b == rs2[9:0]) begin
          coeffs_923 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_924 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h39c == rs2[9:0]) begin
          coeffs_924 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_925 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h39d == rs2[9:0]) begin
          coeffs_925 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_926 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h39e == rs2[9:0]) begin
          coeffs_926 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_927 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h39f == rs2[9:0]) begin
          coeffs_927 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_928 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a0 == rs2[9:0]) begin
          coeffs_928 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_929 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a1 == rs2[9:0]) begin
          coeffs_929 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_930 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a2 == rs2[9:0]) begin
          coeffs_930 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_931 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a3 == rs2[9:0]) begin
          coeffs_931 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_932 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a4 == rs2[9:0]) begin
          coeffs_932 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_933 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a5 == rs2[9:0]) begin
          coeffs_933 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_934 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a6 == rs2[9:0]) begin
          coeffs_934 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_935 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a7 == rs2[9:0]) begin
          coeffs_935 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_936 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a8 == rs2[9:0]) begin
          coeffs_936 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_937 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a9 == rs2[9:0]) begin
          coeffs_937 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_938 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3aa == rs2[9:0]) begin
          coeffs_938 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_939 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3ab == rs2[9:0]) begin
          coeffs_939 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_940 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3ac == rs2[9:0]) begin
          coeffs_940 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_941 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3ad == rs2[9:0]) begin
          coeffs_941 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_942 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3ae == rs2[9:0]) begin
          coeffs_942 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_943 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3af == rs2[9:0]) begin
          coeffs_943 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_944 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b0 == rs2[9:0]) begin
          coeffs_944 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_945 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b1 == rs2[9:0]) begin
          coeffs_945 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_946 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b2 == rs2[9:0]) begin
          coeffs_946 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_947 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b3 == rs2[9:0]) begin
          coeffs_947 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_948 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b4 == rs2[9:0]) begin
          coeffs_948 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_949 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b5 == rs2[9:0]) begin
          coeffs_949 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_950 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b6 == rs2[9:0]) begin
          coeffs_950 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_951 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b7 == rs2[9:0]) begin
          coeffs_951 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_952 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b8 == rs2[9:0]) begin
          coeffs_952 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_953 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b9 == rs2[9:0]) begin
          coeffs_953 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_954 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3ba == rs2[9:0]) begin
          coeffs_954 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_955 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3bb == rs2[9:0]) begin
          coeffs_955 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_956 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3bc == rs2[9:0]) begin
          coeffs_956 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_957 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3bd == rs2[9:0]) begin
          coeffs_957 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_958 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3be == rs2[9:0]) begin
          coeffs_958 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_959 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3bf == rs2[9:0]) begin
          coeffs_959 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_960 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c0 == rs2[9:0]) begin
          coeffs_960 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_961 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c1 == rs2[9:0]) begin
          coeffs_961 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_962 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c2 == rs2[9:0]) begin
          coeffs_962 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_963 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c3 == rs2[9:0]) begin
          coeffs_963 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_964 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c4 == rs2[9:0]) begin
          coeffs_964 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_965 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c5 == rs2[9:0]) begin
          coeffs_965 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_966 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c6 == rs2[9:0]) begin
          coeffs_966 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_967 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c7 == rs2[9:0]) begin
          coeffs_967 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_968 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c8 == rs2[9:0]) begin
          coeffs_968 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_969 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c9 == rs2[9:0]) begin
          coeffs_969 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_970 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3ca == rs2[9:0]) begin
          coeffs_970 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_971 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3cb == rs2[9:0]) begin
          coeffs_971 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_972 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3cc == rs2[9:0]) begin
          coeffs_972 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_973 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3cd == rs2[9:0]) begin
          coeffs_973 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_974 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3ce == rs2[9:0]) begin
          coeffs_974 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_975 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3cf == rs2[9:0]) begin
          coeffs_975 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_976 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d0 == rs2[9:0]) begin
          coeffs_976 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_977 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d1 == rs2[9:0]) begin
          coeffs_977 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_978 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d2 == rs2[9:0]) begin
          coeffs_978 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_979 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d3 == rs2[9:0]) begin
          coeffs_979 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_980 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d4 == rs2[9:0]) begin
          coeffs_980 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_981 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d5 == rs2[9:0]) begin
          coeffs_981 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_982 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d6 == rs2[9:0]) begin
          coeffs_982 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_983 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d7 == rs2[9:0]) begin
          coeffs_983 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_984 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d8 == rs2[9:0]) begin
          coeffs_984 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_985 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d9 == rs2[9:0]) begin
          coeffs_985 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_986 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3da == rs2[9:0]) begin
          coeffs_986 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_987 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3db == rs2[9:0]) begin
          coeffs_987 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_988 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3dc == rs2[9:0]) begin
          coeffs_988 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_989 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3dd == rs2[9:0]) begin
          coeffs_989 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_990 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3de == rs2[9:0]) begin
          coeffs_990 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_991 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3df == rs2[9:0]) begin
          coeffs_991 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_992 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3e0 == rs2[9:0]) begin
          coeffs_992 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_993 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3e1 == rs2[9:0]) begin
          coeffs_993 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_994 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3e2 == rs2[9:0]) begin
          coeffs_994 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_995 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3e3 == rs2[9:0]) begin
          coeffs_995 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_996 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3e4 == rs2[9:0]) begin
          coeffs_996 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_997 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3e5 == rs2[9:0]) begin
          coeffs_997 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_998 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3e6 == rs2[9:0]) begin
          coeffs_998 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_999 <= 32'sh0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3e7 == rs2[9:0]) begin
          coeffs_999 <= rs1;
        end
      end
    end
    if (reset) begin
      data_0 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_0 <= rs1;
        end
      end
    end
    if (reset) begin
      data_1 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_1 <= data_0;
        end
      end
    end
    if (reset) begin
      data_2 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_2 <= data_1;
        end
      end
    end
    if (reset) begin
      data_3 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_3 <= data_2;
        end
      end
    end
    if (reset) begin
      data_4 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_4 <= data_3;
        end
      end
    end
    if (reset) begin
      data_5 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_5 <= data_4;
        end
      end
    end
    if (reset) begin
      data_6 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_6 <= data_5;
        end
      end
    end
    if (reset) begin
      data_7 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_7 <= data_6;
        end
      end
    end
    if (reset) begin
      data_8 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_8 <= data_7;
        end
      end
    end
    if (reset) begin
      data_9 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_9 <= data_8;
        end
      end
    end
    if (reset) begin
      data_10 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_10 <= data_9;
        end
      end
    end
    if (reset) begin
      data_11 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_11 <= data_10;
        end
      end
    end
    if (reset) begin
      data_12 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_12 <= data_11;
        end
      end
    end
    if (reset) begin
      data_13 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_13 <= data_12;
        end
      end
    end
    if (reset) begin
      data_14 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_14 <= data_13;
        end
      end
    end
    if (reset) begin
      data_15 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_15 <= data_14;
        end
      end
    end
    if (reset) begin
      data_16 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_16 <= data_15;
        end
      end
    end
    if (reset) begin
      data_17 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_17 <= data_16;
        end
      end
    end
    if (reset) begin
      data_18 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_18 <= data_17;
        end
      end
    end
    if (reset) begin
      data_19 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_19 <= data_18;
        end
      end
    end
    if (reset) begin
      data_20 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_20 <= data_19;
        end
      end
    end
    if (reset) begin
      data_21 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_21 <= data_20;
        end
      end
    end
    if (reset) begin
      data_22 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_22 <= data_21;
        end
      end
    end
    if (reset) begin
      data_23 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_23 <= data_22;
        end
      end
    end
    if (reset) begin
      data_24 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_24 <= data_23;
        end
      end
    end
    if (reset) begin
      data_25 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_25 <= data_24;
        end
      end
    end
    if (reset) begin
      data_26 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_26 <= data_25;
        end
      end
    end
    if (reset) begin
      data_27 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_27 <= data_26;
        end
      end
    end
    if (reset) begin
      data_28 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_28 <= data_27;
        end
      end
    end
    if (reset) begin
      data_29 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_29 <= data_28;
        end
      end
    end
    if (reset) begin
      data_30 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_30 <= data_29;
        end
      end
    end
    if (reset) begin
      data_31 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_31 <= data_30;
        end
      end
    end
    if (reset) begin
      data_32 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_32 <= data_31;
        end
      end
    end
    if (reset) begin
      data_33 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_33 <= data_32;
        end
      end
    end
    if (reset) begin
      data_34 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_34 <= data_33;
        end
      end
    end
    if (reset) begin
      data_35 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_35 <= data_34;
        end
      end
    end
    if (reset) begin
      data_36 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_36 <= data_35;
        end
      end
    end
    if (reset) begin
      data_37 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_37 <= data_36;
        end
      end
    end
    if (reset) begin
      data_38 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_38 <= data_37;
        end
      end
    end
    if (reset) begin
      data_39 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_39 <= data_38;
        end
      end
    end
    if (reset) begin
      data_40 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_40 <= data_39;
        end
      end
    end
    if (reset) begin
      data_41 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_41 <= data_40;
        end
      end
    end
    if (reset) begin
      data_42 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_42 <= data_41;
        end
      end
    end
    if (reset) begin
      data_43 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_43 <= data_42;
        end
      end
    end
    if (reset) begin
      data_44 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_44 <= data_43;
        end
      end
    end
    if (reset) begin
      data_45 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_45 <= data_44;
        end
      end
    end
    if (reset) begin
      data_46 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_46 <= data_45;
        end
      end
    end
    if (reset) begin
      data_47 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_47 <= data_46;
        end
      end
    end
    if (reset) begin
      data_48 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_48 <= data_47;
        end
      end
    end
    if (reset) begin
      data_49 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_49 <= data_48;
        end
      end
    end
    if (reset) begin
      data_50 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_50 <= data_49;
        end
      end
    end
    if (reset) begin
      data_51 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_51 <= data_50;
        end
      end
    end
    if (reset) begin
      data_52 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_52 <= data_51;
        end
      end
    end
    if (reset) begin
      data_53 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_53 <= data_52;
        end
      end
    end
    if (reset) begin
      data_54 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_54 <= data_53;
        end
      end
    end
    if (reset) begin
      data_55 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_55 <= data_54;
        end
      end
    end
    if (reset) begin
      data_56 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_56 <= data_55;
        end
      end
    end
    if (reset) begin
      data_57 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_57 <= data_56;
        end
      end
    end
    if (reset) begin
      data_58 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_58 <= data_57;
        end
      end
    end
    if (reset) begin
      data_59 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_59 <= data_58;
        end
      end
    end
    if (reset) begin
      data_60 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_60 <= data_59;
        end
      end
    end
    if (reset) begin
      data_61 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_61 <= data_60;
        end
      end
    end
    if (reset) begin
      data_62 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_62 <= data_61;
        end
      end
    end
    if (reset) begin
      data_63 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_63 <= data_62;
        end
      end
    end
    if (reset) begin
      data_64 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_64 <= data_63;
        end
      end
    end
    if (reset) begin
      data_65 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_65 <= data_64;
        end
      end
    end
    if (reset) begin
      data_66 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_66 <= data_65;
        end
      end
    end
    if (reset) begin
      data_67 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_67 <= data_66;
        end
      end
    end
    if (reset) begin
      data_68 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_68 <= data_67;
        end
      end
    end
    if (reset) begin
      data_69 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_69 <= data_68;
        end
      end
    end
    if (reset) begin
      data_70 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_70 <= data_69;
        end
      end
    end
    if (reset) begin
      data_71 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_71 <= data_70;
        end
      end
    end
    if (reset) begin
      data_72 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_72 <= data_71;
        end
      end
    end
    if (reset) begin
      data_73 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_73 <= data_72;
        end
      end
    end
    if (reset) begin
      data_74 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_74 <= data_73;
        end
      end
    end
    if (reset) begin
      data_75 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_75 <= data_74;
        end
      end
    end
    if (reset) begin
      data_76 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_76 <= data_75;
        end
      end
    end
    if (reset) begin
      data_77 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_77 <= data_76;
        end
      end
    end
    if (reset) begin
      data_78 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_78 <= data_77;
        end
      end
    end
    if (reset) begin
      data_79 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_79 <= data_78;
        end
      end
    end
    if (reset) begin
      data_80 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_80 <= data_79;
        end
      end
    end
    if (reset) begin
      data_81 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_81 <= data_80;
        end
      end
    end
    if (reset) begin
      data_82 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_82 <= data_81;
        end
      end
    end
    if (reset) begin
      data_83 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_83 <= data_82;
        end
      end
    end
    if (reset) begin
      data_84 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_84 <= data_83;
        end
      end
    end
    if (reset) begin
      data_85 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_85 <= data_84;
        end
      end
    end
    if (reset) begin
      data_86 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_86 <= data_85;
        end
      end
    end
    if (reset) begin
      data_87 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_87 <= data_86;
        end
      end
    end
    if (reset) begin
      data_88 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_88 <= data_87;
        end
      end
    end
    if (reset) begin
      data_89 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_89 <= data_88;
        end
      end
    end
    if (reset) begin
      data_90 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_90 <= data_89;
        end
      end
    end
    if (reset) begin
      data_91 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_91 <= data_90;
        end
      end
    end
    if (reset) begin
      data_92 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_92 <= data_91;
        end
      end
    end
    if (reset) begin
      data_93 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_93 <= data_92;
        end
      end
    end
    if (reset) begin
      data_94 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_94 <= data_93;
        end
      end
    end
    if (reset) begin
      data_95 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_95 <= data_94;
        end
      end
    end
    if (reset) begin
      data_96 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_96 <= data_95;
        end
      end
    end
    if (reset) begin
      data_97 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_97 <= data_96;
        end
      end
    end
    if (reset) begin
      data_98 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_98 <= data_97;
        end
      end
    end
    if (reset) begin
      data_99 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_99 <= data_98;
        end
      end
    end
    if (reset) begin
      data_100 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_100 <= data_99;
        end
      end
    end
    if (reset) begin
      data_101 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_101 <= data_100;
        end
      end
    end
    if (reset) begin
      data_102 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_102 <= data_101;
        end
      end
    end
    if (reset) begin
      data_103 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_103 <= data_102;
        end
      end
    end
    if (reset) begin
      data_104 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_104 <= data_103;
        end
      end
    end
    if (reset) begin
      data_105 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_105 <= data_104;
        end
      end
    end
    if (reset) begin
      data_106 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_106 <= data_105;
        end
      end
    end
    if (reset) begin
      data_107 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_107 <= data_106;
        end
      end
    end
    if (reset) begin
      data_108 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_108 <= data_107;
        end
      end
    end
    if (reset) begin
      data_109 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_109 <= data_108;
        end
      end
    end
    if (reset) begin
      data_110 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_110 <= data_109;
        end
      end
    end
    if (reset) begin
      data_111 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_111 <= data_110;
        end
      end
    end
    if (reset) begin
      data_112 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_112 <= data_111;
        end
      end
    end
    if (reset) begin
      data_113 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_113 <= data_112;
        end
      end
    end
    if (reset) begin
      data_114 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_114 <= data_113;
        end
      end
    end
    if (reset) begin
      data_115 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_115 <= data_114;
        end
      end
    end
    if (reset) begin
      data_116 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_116 <= data_115;
        end
      end
    end
    if (reset) begin
      data_117 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_117 <= data_116;
        end
      end
    end
    if (reset) begin
      data_118 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_118 <= data_117;
        end
      end
    end
    if (reset) begin
      data_119 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_119 <= data_118;
        end
      end
    end
    if (reset) begin
      data_120 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_120 <= data_119;
        end
      end
    end
    if (reset) begin
      data_121 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_121 <= data_120;
        end
      end
    end
    if (reset) begin
      data_122 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_122 <= data_121;
        end
      end
    end
    if (reset) begin
      data_123 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_123 <= data_122;
        end
      end
    end
    if (reset) begin
      data_124 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_124 <= data_123;
        end
      end
    end
    if (reset) begin
      data_125 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_125 <= data_124;
        end
      end
    end
    if (reset) begin
      data_126 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_126 <= data_125;
        end
      end
    end
    if (reset) begin
      data_127 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_127 <= data_126;
        end
      end
    end
    if (reset) begin
      data_128 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_128 <= data_127;
        end
      end
    end
    if (reset) begin
      data_129 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_129 <= data_128;
        end
      end
    end
    if (reset) begin
      data_130 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_130 <= data_129;
        end
      end
    end
    if (reset) begin
      data_131 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_131 <= data_130;
        end
      end
    end
    if (reset) begin
      data_132 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_132 <= data_131;
        end
      end
    end
    if (reset) begin
      data_133 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_133 <= data_132;
        end
      end
    end
    if (reset) begin
      data_134 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_134 <= data_133;
        end
      end
    end
    if (reset) begin
      data_135 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_135 <= data_134;
        end
      end
    end
    if (reset) begin
      data_136 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_136 <= data_135;
        end
      end
    end
    if (reset) begin
      data_137 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_137 <= data_136;
        end
      end
    end
    if (reset) begin
      data_138 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_138 <= data_137;
        end
      end
    end
    if (reset) begin
      data_139 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_139 <= data_138;
        end
      end
    end
    if (reset) begin
      data_140 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_140 <= data_139;
        end
      end
    end
    if (reset) begin
      data_141 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_141 <= data_140;
        end
      end
    end
    if (reset) begin
      data_142 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_142 <= data_141;
        end
      end
    end
    if (reset) begin
      data_143 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_143 <= data_142;
        end
      end
    end
    if (reset) begin
      data_144 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_144 <= data_143;
        end
      end
    end
    if (reset) begin
      data_145 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_145 <= data_144;
        end
      end
    end
    if (reset) begin
      data_146 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_146 <= data_145;
        end
      end
    end
    if (reset) begin
      data_147 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_147 <= data_146;
        end
      end
    end
    if (reset) begin
      data_148 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_148 <= data_147;
        end
      end
    end
    if (reset) begin
      data_149 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_149 <= data_148;
        end
      end
    end
    if (reset) begin
      data_150 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_150 <= data_149;
        end
      end
    end
    if (reset) begin
      data_151 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_151 <= data_150;
        end
      end
    end
    if (reset) begin
      data_152 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_152 <= data_151;
        end
      end
    end
    if (reset) begin
      data_153 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_153 <= data_152;
        end
      end
    end
    if (reset) begin
      data_154 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_154 <= data_153;
        end
      end
    end
    if (reset) begin
      data_155 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_155 <= data_154;
        end
      end
    end
    if (reset) begin
      data_156 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_156 <= data_155;
        end
      end
    end
    if (reset) begin
      data_157 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_157 <= data_156;
        end
      end
    end
    if (reset) begin
      data_158 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_158 <= data_157;
        end
      end
    end
    if (reset) begin
      data_159 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_159 <= data_158;
        end
      end
    end
    if (reset) begin
      data_160 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_160 <= data_159;
        end
      end
    end
    if (reset) begin
      data_161 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_161 <= data_160;
        end
      end
    end
    if (reset) begin
      data_162 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_162 <= data_161;
        end
      end
    end
    if (reset) begin
      data_163 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_163 <= data_162;
        end
      end
    end
    if (reset) begin
      data_164 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_164 <= data_163;
        end
      end
    end
    if (reset) begin
      data_165 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_165 <= data_164;
        end
      end
    end
    if (reset) begin
      data_166 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_166 <= data_165;
        end
      end
    end
    if (reset) begin
      data_167 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_167 <= data_166;
        end
      end
    end
    if (reset) begin
      data_168 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_168 <= data_167;
        end
      end
    end
    if (reset) begin
      data_169 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_169 <= data_168;
        end
      end
    end
    if (reset) begin
      data_170 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_170 <= data_169;
        end
      end
    end
    if (reset) begin
      data_171 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_171 <= data_170;
        end
      end
    end
    if (reset) begin
      data_172 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_172 <= data_171;
        end
      end
    end
    if (reset) begin
      data_173 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_173 <= data_172;
        end
      end
    end
    if (reset) begin
      data_174 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_174 <= data_173;
        end
      end
    end
    if (reset) begin
      data_175 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_175 <= data_174;
        end
      end
    end
    if (reset) begin
      data_176 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_176 <= data_175;
        end
      end
    end
    if (reset) begin
      data_177 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_177 <= data_176;
        end
      end
    end
    if (reset) begin
      data_178 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_178 <= data_177;
        end
      end
    end
    if (reset) begin
      data_179 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_179 <= data_178;
        end
      end
    end
    if (reset) begin
      data_180 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_180 <= data_179;
        end
      end
    end
    if (reset) begin
      data_181 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_181 <= data_180;
        end
      end
    end
    if (reset) begin
      data_182 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_182 <= data_181;
        end
      end
    end
    if (reset) begin
      data_183 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_183 <= data_182;
        end
      end
    end
    if (reset) begin
      data_184 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_184 <= data_183;
        end
      end
    end
    if (reset) begin
      data_185 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_185 <= data_184;
        end
      end
    end
    if (reset) begin
      data_186 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_186 <= data_185;
        end
      end
    end
    if (reset) begin
      data_187 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_187 <= data_186;
        end
      end
    end
    if (reset) begin
      data_188 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_188 <= data_187;
        end
      end
    end
    if (reset) begin
      data_189 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_189 <= data_188;
        end
      end
    end
    if (reset) begin
      data_190 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_190 <= data_189;
        end
      end
    end
    if (reset) begin
      data_191 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_191 <= data_190;
        end
      end
    end
    if (reset) begin
      data_192 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_192 <= data_191;
        end
      end
    end
    if (reset) begin
      data_193 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_193 <= data_192;
        end
      end
    end
    if (reset) begin
      data_194 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_194 <= data_193;
        end
      end
    end
    if (reset) begin
      data_195 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_195 <= data_194;
        end
      end
    end
    if (reset) begin
      data_196 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_196 <= data_195;
        end
      end
    end
    if (reset) begin
      data_197 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_197 <= data_196;
        end
      end
    end
    if (reset) begin
      data_198 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_198 <= data_197;
        end
      end
    end
    if (reset) begin
      data_199 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_199 <= data_198;
        end
      end
    end
    if (reset) begin
      data_200 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_200 <= data_199;
        end
      end
    end
    if (reset) begin
      data_201 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_201 <= data_200;
        end
      end
    end
    if (reset) begin
      data_202 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_202 <= data_201;
        end
      end
    end
    if (reset) begin
      data_203 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_203 <= data_202;
        end
      end
    end
    if (reset) begin
      data_204 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_204 <= data_203;
        end
      end
    end
    if (reset) begin
      data_205 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_205 <= data_204;
        end
      end
    end
    if (reset) begin
      data_206 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_206 <= data_205;
        end
      end
    end
    if (reset) begin
      data_207 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_207 <= data_206;
        end
      end
    end
    if (reset) begin
      data_208 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_208 <= data_207;
        end
      end
    end
    if (reset) begin
      data_209 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_209 <= data_208;
        end
      end
    end
    if (reset) begin
      data_210 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_210 <= data_209;
        end
      end
    end
    if (reset) begin
      data_211 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_211 <= data_210;
        end
      end
    end
    if (reset) begin
      data_212 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_212 <= data_211;
        end
      end
    end
    if (reset) begin
      data_213 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_213 <= data_212;
        end
      end
    end
    if (reset) begin
      data_214 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_214 <= data_213;
        end
      end
    end
    if (reset) begin
      data_215 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_215 <= data_214;
        end
      end
    end
    if (reset) begin
      data_216 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_216 <= data_215;
        end
      end
    end
    if (reset) begin
      data_217 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_217 <= data_216;
        end
      end
    end
    if (reset) begin
      data_218 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_218 <= data_217;
        end
      end
    end
    if (reset) begin
      data_219 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_219 <= data_218;
        end
      end
    end
    if (reset) begin
      data_220 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_220 <= data_219;
        end
      end
    end
    if (reset) begin
      data_221 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_221 <= data_220;
        end
      end
    end
    if (reset) begin
      data_222 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_222 <= data_221;
        end
      end
    end
    if (reset) begin
      data_223 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_223 <= data_222;
        end
      end
    end
    if (reset) begin
      data_224 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_224 <= data_223;
        end
      end
    end
    if (reset) begin
      data_225 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_225 <= data_224;
        end
      end
    end
    if (reset) begin
      data_226 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_226 <= data_225;
        end
      end
    end
    if (reset) begin
      data_227 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_227 <= data_226;
        end
      end
    end
    if (reset) begin
      data_228 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_228 <= data_227;
        end
      end
    end
    if (reset) begin
      data_229 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_229 <= data_228;
        end
      end
    end
    if (reset) begin
      data_230 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_230 <= data_229;
        end
      end
    end
    if (reset) begin
      data_231 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_231 <= data_230;
        end
      end
    end
    if (reset) begin
      data_232 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_232 <= data_231;
        end
      end
    end
    if (reset) begin
      data_233 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_233 <= data_232;
        end
      end
    end
    if (reset) begin
      data_234 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_234 <= data_233;
        end
      end
    end
    if (reset) begin
      data_235 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_235 <= data_234;
        end
      end
    end
    if (reset) begin
      data_236 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_236 <= data_235;
        end
      end
    end
    if (reset) begin
      data_237 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_237 <= data_236;
        end
      end
    end
    if (reset) begin
      data_238 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_238 <= data_237;
        end
      end
    end
    if (reset) begin
      data_239 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_239 <= data_238;
        end
      end
    end
    if (reset) begin
      data_240 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_240 <= data_239;
        end
      end
    end
    if (reset) begin
      data_241 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_241 <= data_240;
        end
      end
    end
    if (reset) begin
      data_242 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_242 <= data_241;
        end
      end
    end
    if (reset) begin
      data_243 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_243 <= data_242;
        end
      end
    end
    if (reset) begin
      data_244 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_244 <= data_243;
        end
      end
    end
    if (reset) begin
      data_245 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_245 <= data_244;
        end
      end
    end
    if (reset) begin
      data_246 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_246 <= data_245;
        end
      end
    end
    if (reset) begin
      data_247 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_247 <= data_246;
        end
      end
    end
    if (reset) begin
      data_248 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_248 <= data_247;
        end
      end
    end
    if (reset) begin
      data_249 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_249 <= data_248;
        end
      end
    end
    if (reset) begin
      data_250 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_250 <= data_249;
        end
      end
    end
    if (reset) begin
      data_251 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_251 <= data_250;
        end
      end
    end
    if (reset) begin
      data_252 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_252 <= data_251;
        end
      end
    end
    if (reset) begin
      data_253 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_253 <= data_252;
        end
      end
    end
    if (reset) begin
      data_254 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_254 <= data_253;
        end
      end
    end
    if (reset) begin
      data_255 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_255 <= data_254;
        end
      end
    end
    if (reset) begin
      data_256 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_256 <= data_255;
        end
      end
    end
    if (reset) begin
      data_257 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_257 <= data_256;
        end
      end
    end
    if (reset) begin
      data_258 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_258 <= data_257;
        end
      end
    end
    if (reset) begin
      data_259 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_259 <= data_258;
        end
      end
    end
    if (reset) begin
      data_260 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_260 <= data_259;
        end
      end
    end
    if (reset) begin
      data_261 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_261 <= data_260;
        end
      end
    end
    if (reset) begin
      data_262 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_262 <= data_261;
        end
      end
    end
    if (reset) begin
      data_263 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_263 <= data_262;
        end
      end
    end
    if (reset) begin
      data_264 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_264 <= data_263;
        end
      end
    end
    if (reset) begin
      data_265 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_265 <= data_264;
        end
      end
    end
    if (reset) begin
      data_266 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_266 <= data_265;
        end
      end
    end
    if (reset) begin
      data_267 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_267 <= data_266;
        end
      end
    end
    if (reset) begin
      data_268 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_268 <= data_267;
        end
      end
    end
    if (reset) begin
      data_269 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_269 <= data_268;
        end
      end
    end
    if (reset) begin
      data_270 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_270 <= data_269;
        end
      end
    end
    if (reset) begin
      data_271 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_271 <= data_270;
        end
      end
    end
    if (reset) begin
      data_272 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_272 <= data_271;
        end
      end
    end
    if (reset) begin
      data_273 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_273 <= data_272;
        end
      end
    end
    if (reset) begin
      data_274 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_274 <= data_273;
        end
      end
    end
    if (reset) begin
      data_275 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_275 <= data_274;
        end
      end
    end
    if (reset) begin
      data_276 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_276 <= data_275;
        end
      end
    end
    if (reset) begin
      data_277 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_277 <= data_276;
        end
      end
    end
    if (reset) begin
      data_278 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_278 <= data_277;
        end
      end
    end
    if (reset) begin
      data_279 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_279 <= data_278;
        end
      end
    end
    if (reset) begin
      data_280 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_280 <= data_279;
        end
      end
    end
    if (reset) begin
      data_281 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_281 <= data_280;
        end
      end
    end
    if (reset) begin
      data_282 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_282 <= data_281;
        end
      end
    end
    if (reset) begin
      data_283 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_283 <= data_282;
        end
      end
    end
    if (reset) begin
      data_284 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_284 <= data_283;
        end
      end
    end
    if (reset) begin
      data_285 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_285 <= data_284;
        end
      end
    end
    if (reset) begin
      data_286 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_286 <= data_285;
        end
      end
    end
    if (reset) begin
      data_287 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_287 <= data_286;
        end
      end
    end
    if (reset) begin
      data_288 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_288 <= data_287;
        end
      end
    end
    if (reset) begin
      data_289 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_289 <= data_288;
        end
      end
    end
    if (reset) begin
      data_290 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_290 <= data_289;
        end
      end
    end
    if (reset) begin
      data_291 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_291 <= data_290;
        end
      end
    end
    if (reset) begin
      data_292 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_292 <= data_291;
        end
      end
    end
    if (reset) begin
      data_293 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_293 <= data_292;
        end
      end
    end
    if (reset) begin
      data_294 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_294 <= data_293;
        end
      end
    end
    if (reset) begin
      data_295 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_295 <= data_294;
        end
      end
    end
    if (reset) begin
      data_296 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_296 <= data_295;
        end
      end
    end
    if (reset) begin
      data_297 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_297 <= data_296;
        end
      end
    end
    if (reset) begin
      data_298 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_298 <= data_297;
        end
      end
    end
    if (reset) begin
      data_299 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_299 <= data_298;
        end
      end
    end
    if (reset) begin
      data_300 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_300 <= data_299;
        end
      end
    end
    if (reset) begin
      data_301 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_301 <= data_300;
        end
      end
    end
    if (reset) begin
      data_302 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_302 <= data_301;
        end
      end
    end
    if (reset) begin
      data_303 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_303 <= data_302;
        end
      end
    end
    if (reset) begin
      data_304 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_304 <= data_303;
        end
      end
    end
    if (reset) begin
      data_305 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_305 <= data_304;
        end
      end
    end
    if (reset) begin
      data_306 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_306 <= data_305;
        end
      end
    end
    if (reset) begin
      data_307 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_307 <= data_306;
        end
      end
    end
    if (reset) begin
      data_308 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_308 <= data_307;
        end
      end
    end
    if (reset) begin
      data_309 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_309 <= data_308;
        end
      end
    end
    if (reset) begin
      data_310 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_310 <= data_309;
        end
      end
    end
    if (reset) begin
      data_311 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_311 <= data_310;
        end
      end
    end
    if (reset) begin
      data_312 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_312 <= data_311;
        end
      end
    end
    if (reset) begin
      data_313 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_313 <= data_312;
        end
      end
    end
    if (reset) begin
      data_314 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_314 <= data_313;
        end
      end
    end
    if (reset) begin
      data_315 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_315 <= data_314;
        end
      end
    end
    if (reset) begin
      data_316 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_316 <= data_315;
        end
      end
    end
    if (reset) begin
      data_317 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_317 <= data_316;
        end
      end
    end
    if (reset) begin
      data_318 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_318 <= data_317;
        end
      end
    end
    if (reset) begin
      data_319 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_319 <= data_318;
        end
      end
    end
    if (reset) begin
      data_320 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_320 <= data_319;
        end
      end
    end
    if (reset) begin
      data_321 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_321 <= data_320;
        end
      end
    end
    if (reset) begin
      data_322 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_322 <= data_321;
        end
      end
    end
    if (reset) begin
      data_323 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_323 <= data_322;
        end
      end
    end
    if (reset) begin
      data_324 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_324 <= data_323;
        end
      end
    end
    if (reset) begin
      data_325 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_325 <= data_324;
        end
      end
    end
    if (reset) begin
      data_326 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_326 <= data_325;
        end
      end
    end
    if (reset) begin
      data_327 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_327 <= data_326;
        end
      end
    end
    if (reset) begin
      data_328 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_328 <= data_327;
        end
      end
    end
    if (reset) begin
      data_329 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_329 <= data_328;
        end
      end
    end
    if (reset) begin
      data_330 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_330 <= data_329;
        end
      end
    end
    if (reset) begin
      data_331 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_331 <= data_330;
        end
      end
    end
    if (reset) begin
      data_332 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_332 <= data_331;
        end
      end
    end
    if (reset) begin
      data_333 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_333 <= data_332;
        end
      end
    end
    if (reset) begin
      data_334 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_334 <= data_333;
        end
      end
    end
    if (reset) begin
      data_335 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_335 <= data_334;
        end
      end
    end
    if (reset) begin
      data_336 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_336 <= data_335;
        end
      end
    end
    if (reset) begin
      data_337 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_337 <= data_336;
        end
      end
    end
    if (reset) begin
      data_338 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_338 <= data_337;
        end
      end
    end
    if (reset) begin
      data_339 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_339 <= data_338;
        end
      end
    end
    if (reset) begin
      data_340 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_340 <= data_339;
        end
      end
    end
    if (reset) begin
      data_341 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_341 <= data_340;
        end
      end
    end
    if (reset) begin
      data_342 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_342 <= data_341;
        end
      end
    end
    if (reset) begin
      data_343 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_343 <= data_342;
        end
      end
    end
    if (reset) begin
      data_344 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_344 <= data_343;
        end
      end
    end
    if (reset) begin
      data_345 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_345 <= data_344;
        end
      end
    end
    if (reset) begin
      data_346 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_346 <= data_345;
        end
      end
    end
    if (reset) begin
      data_347 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_347 <= data_346;
        end
      end
    end
    if (reset) begin
      data_348 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_348 <= data_347;
        end
      end
    end
    if (reset) begin
      data_349 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_349 <= data_348;
        end
      end
    end
    if (reset) begin
      data_350 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_350 <= data_349;
        end
      end
    end
    if (reset) begin
      data_351 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_351 <= data_350;
        end
      end
    end
    if (reset) begin
      data_352 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_352 <= data_351;
        end
      end
    end
    if (reset) begin
      data_353 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_353 <= data_352;
        end
      end
    end
    if (reset) begin
      data_354 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_354 <= data_353;
        end
      end
    end
    if (reset) begin
      data_355 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_355 <= data_354;
        end
      end
    end
    if (reset) begin
      data_356 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_356 <= data_355;
        end
      end
    end
    if (reset) begin
      data_357 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_357 <= data_356;
        end
      end
    end
    if (reset) begin
      data_358 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_358 <= data_357;
        end
      end
    end
    if (reset) begin
      data_359 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_359 <= data_358;
        end
      end
    end
    if (reset) begin
      data_360 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_360 <= data_359;
        end
      end
    end
    if (reset) begin
      data_361 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_361 <= data_360;
        end
      end
    end
    if (reset) begin
      data_362 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_362 <= data_361;
        end
      end
    end
    if (reset) begin
      data_363 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_363 <= data_362;
        end
      end
    end
    if (reset) begin
      data_364 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_364 <= data_363;
        end
      end
    end
    if (reset) begin
      data_365 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_365 <= data_364;
        end
      end
    end
    if (reset) begin
      data_366 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_366 <= data_365;
        end
      end
    end
    if (reset) begin
      data_367 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_367 <= data_366;
        end
      end
    end
    if (reset) begin
      data_368 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_368 <= data_367;
        end
      end
    end
    if (reset) begin
      data_369 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_369 <= data_368;
        end
      end
    end
    if (reset) begin
      data_370 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_370 <= data_369;
        end
      end
    end
    if (reset) begin
      data_371 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_371 <= data_370;
        end
      end
    end
    if (reset) begin
      data_372 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_372 <= data_371;
        end
      end
    end
    if (reset) begin
      data_373 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_373 <= data_372;
        end
      end
    end
    if (reset) begin
      data_374 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_374 <= data_373;
        end
      end
    end
    if (reset) begin
      data_375 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_375 <= data_374;
        end
      end
    end
    if (reset) begin
      data_376 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_376 <= data_375;
        end
      end
    end
    if (reset) begin
      data_377 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_377 <= data_376;
        end
      end
    end
    if (reset) begin
      data_378 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_378 <= data_377;
        end
      end
    end
    if (reset) begin
      data_379 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_379 <= data_378;
        end
      end
    end
    if (reset) begin
      data_380 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_380 <= data_379;
        end
      end
    end
    if (reset) begin
      data_381 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_381 <= data_380;
        end
      end
    end
    if (reset) begin
      data_382 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_382 <= data_381;
        end
      end
    end
    if (reset) begin
      data_383 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_383 <= data_382;
        end
      end
    end
    if (reset) begin
      data_384 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_384 <= data_383;
        end
      end
    end
    if (reset) begin
      data_385 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_385 <= data_384;
        end
      end
    end
    if (reset) begin
      data_386 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_386 <= data_385;
        end
      end
    end
    if (reset) begin
      data_387 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_387 <= data_386;
        end
      end
    end
    if (reset) begin
      data_388 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_388 <= data_387;
        end
      end
    end
    if (reset) begin
      data_389 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_389 <= data_388;
        end
      end
    end
    if (reset) begin
      data_390 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_390 <= data_389;
        end
      end
    end
    if (reset) begin
      data_391 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_391 <= data_390;
        end
      end
    end
    if (reset) begin
      data_392 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_392 <= data_391;
        end
      end
    end
    if (reset) begin
      data_393 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_393 <= data_392;
        end
      end
    end
    if (reset) begin
      data_394 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_394 <= data_393;
        end
      end
    end
    if (reset) begin
      data_395 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_395 <= data_394;
        end
      end
    end
    if (reset) begin
      data_396 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_396 <= data_395;
        end
      end
    end
    if (reset) begin
      data_397 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_397 <= data_396;
        end
      end
    end
    if (reset) begin
      data_398 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_398 <= data_397;
        end
      end
    end
    if (reset) begin
      data_399 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_399 <= data_398;
        end
      end
    end
    if (reset) begin
      data_400 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_400 <= data_399;
        end
      end
    end
    if (reset) begin
      data_401 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_401 <= data_400;
        end
      end
    end
    if (reset) begin
      data_402 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_402 <= data_401;
        end
      end
    end
    if (reset) begin
      data_403 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_403 <= data_402;
        end
      end
    end
    if (reset) begin
      data_404 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_404 <= data_403;
        end
      end
    end
    if (reset) begin
      data_405 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_405 <= data_404;
        end
      end
    end
    if (reset) begin
      data_406 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_406 <= data_405;
        end
      end
    end
    if (reset) begin
      data_407 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_407 <= data_406;
        end
      end
    end
    if (reset) begin
      data_408 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_408 <= data_407;
        end
      end
    end
    if (reset) begin
      data_409 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_409 <= data_408;
        end
      end
    end
    if (reset) begin
      data_410 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_410 <= data_409;
        end
      end
    end
    if (reset) begin
      data_411 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_411 <= data_410;
        end
      end
    end
    if (reset) begin
      data_412 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_412 <= data_411;
        end
      end
    end
    if (reset) begin
      data_413 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_413 <= data_412;
        end
      end
    end
    if (reset) begin
      data_414 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_414 <= data_413;
        end
      end
    end
    if (reset) begin
      data_415 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_415 <= data_414;
        end
      end
    end
    if (reset) begin
      data_416 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_416 <= data_415;
        end
      end
    end
    if (reset) begin
      data_417 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_417 <= data_416;
        end
      end
    end
    if (reset) begin
      data_418 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_418 <= data_417;
        end
      end
    end
    if (reset) begin
      data_419 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_419 <= data_418;
        end
      end
    end
    if (reset) begin
      data_420 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_420 <= data_419;
        end
      end
    end
    if (reset) begin
      data_421 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_421 <= data_420;
        end
      end
    end
    if (reset) begin
      data_422 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_422 <= data_421;
        end
      end
    end
    if (reset) begin
      data_423 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_423 <= data_422;
        end
      end
    end
    if (reset) begin
      data_424 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_424 <= data_423;
        end
      end
    end
    if (reset) begin
      data_425 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_425 <= data_424;
        end
      end
    end
    if (reset) begin
      data_426 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_426 <= data_425;
        end
      end
    end
    if (reset) begin
      data_427 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_427 <= data_426;
        end
      end
    end
    if (reset) begin
      data_428 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_428 <= data_427;
        end
      end
    end
    if (reset) begin
      data_429 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_429 <= data_428;
        end
      end
    end
    if (reset) begin
      data_430 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_430 <= data_429;
        end
      end
    end
    if (reset) begin
      data_431 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_431 <= data_430;
        end
      end
    end
    if (reset) begin
      data_432 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_432 <= data_431;
        end
      end
    end
    if (reset) begin
      data_433 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_433 <= data_432;
        end
      end
    end
    if (reset) begin
      data_434 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_434 <= data_433;
        end
      end
    end
    if (reset) begin
      data_435 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_435 <= data_434;
        end
      end
    end
    if (reset) begin
      data_436 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_436 <= data_435;
        end
      end
    end
    if (reset) begin
      data_437 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_437 <= data_436;
        end
      end
    end
    if (reset) begin
      data_438 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_438 <= data_437;
        end
      end
    end
    if (reset) begin
      data_439 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_439 <= data_438;
        end
      end
    end
    if (reset) begin
      data_440 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_440 <= data_439;
        end
      end
    end
    if (reset) begin
      data_441 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_441 <= data_440;
        end
      end
    end
    if (reset) begin
      data_442 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_442 <= data_441;
        end
      end
    end
    if (reset) begin
      data_443 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_443 <= data_442;
        end
      end
    end
    if (reset) begin
      data_444 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_444 <= data_443;
        end
      end
    end
    if (reset) begin
      data_445 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_445 <= data_444;
        end
      end
    end
    if (reset) begin
      data_446 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_446 <= data_445;
        end
      end
    end
    if (reset) begin
      data_447 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_447 <= data_446;
        end
      end
    end
    if (reset) begin
      data_448 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_448 <= data_447;
        end
      end
    end
    if (reset) begin
      data_449 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_449 <= data_448;
        end
      end
    end
    if (reset) begin
      data_450 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_450 <= data_449;
        end
      end
    end
    if (reset) begin
      data_451 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_451 <= data_450;
        end
      end
    end
    if (reset) begin
      data_452 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_452 <= data_451;
        end
      end
    end
    if (reset) begin
      data_453 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_453 <= data_452;
        end
      end
    end
    if (reset) begin
      data_454 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_454 <= data_453;
        end
      end
    end
    if (reset) begin
      data_455 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_455 <= data_454;
        end
      end
    end
    if (reset) begin
      data_456 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_456 <= data_455;
        end
      end
    end
    if (reset) begin
      data_457 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_457 <= data_456;
        end
      end
    end
    if (reset) begin
      data_458 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_458 <= data_457;
        end
      end
    end
    if (reset) begin
      data_459 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_459 <= data_458;
        end
      end
    end
    if (reset) begin
      data_460 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_460 <= data_459;
        end
      end
    end
    if (reset) begin
      data_461 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_461 <= data_460;
        end
      end
    end
    if (reset) begin
      data_462 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_462 <= data_461;
        end
      end
    end
    if (reset) begin
      data_463 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_463 <= data_462;
        end
      end
    end
    if (reset) begin
      data_464 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_464 <= data_463;
        end
      end
    end
    if (reset) begin
      data_465 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_465 <= data_464;
        end
      end
    end
    if (reset) begin
      data_466 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_466 <= data_465;
        end
      end
    end
    if (reset) begin
      data_467 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_467 <= data_466;
        end
      end
    end
    if (reset) begin
      data_468 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_468 <= data_467;
        end
      end
    end
    if (reset) begin
      data_469 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_469 <= data_468;
        end
      end
    end
    if (reset) begin
      data_470 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_470 <= data_469;
        end
      end
    end
    if (reset) begin
      data_471 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_471 <= data_470;
        end
      end
    end
    if (reset) begin
      data_472 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_472 <= data_471;
        end
      end
    end
    if (reset) begin
      data_473 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_473 <= data_472;
        end
      end
    end
    if (reset) begin
      data_474 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_474 <= data_473;
        end
      end
    end
    if (reset) begin
      data_475 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_475 <= data_474;
        end
      end
    end
    if (reset) begin
      data_476 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_476 <= data_475;
        end
      end
    end
    if (reset) begin
      data_477 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_477 <= data_476;
        end
      end
    end
    if (reset) begin
      data_478 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_478 <= data_477;
        end
      end
    end
    if (reset) begin
      data_479 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_479 <= data_478;
        end
      end
    end
    if (reset) begin
      data_480 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_480 <= data_479;
        end
      end
    end
    if (reset) begin
      data_481 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_481 <= data_480;
        end
      end
    end
    if (reset) begin
      data_482 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_482 <= data_481;
        end
      end
    end
    if (reset) begin
      data_483 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_483 <= data_482;
        end
      end
    end
    if (reset) begin
      data_484 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_484 <= data_483;
        end
      end
    end
    if (reset) begin
      data_485 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_485 <= data_484;
        end
      end
    end
    if (reset) begin
      data_486 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_486 <= data_485;
        end
      end
    end
    if (reset) begin
      data_487 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_487 <= data_486;
        end
      end
    end
    if (reset) begin
      data_488 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_488 <= data_487;
        end
      end
    end
    if (reset) begin
      data_489 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_489 <= data_488;
        end
      end
    end
    if (reset) begin
      data_490 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_490 <= data_489;
        end
      end
    end
    if (reset) begin
      data_491 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_491 <= data_490;
        end
      end
    end
    if (reset) begin
      data_492 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_492 <= data_491;
        end
      end
    end
    if (reset) begin
      data_493 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_493 <= data_492;
        end
      end
    end
    if (reset) begin
      data_494 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_494 <= data_493;
        end
      end
    end
    if (reset) begin
      data_495 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_495 <= data_494;
        end
      end
    end
    if (reset) begin
      data_496 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_496 <= data_495;
        end
      end
    end
    if (reset) begin
      data_497 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_497 <= data_496;
        end
      end
    end
    if (reset) begin
      data_498 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_498 <= data_497;
        end
      end
    end
    if (reset) begin
      data_499 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_499 <= data_498;
        end
      end
    end
    if (reset) begin
      data_500 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_500 <= data_499;
        end
      end
    end
    if (reset) begin
      data_501 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_501 <= data_500;
        end
      end
    end
    if (reset) begin
      data_502 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_502 <= data_501;
        end
      end
    end
    if (reset) begin
      data_503 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_503 <= data_502;
        end
      end
    end
    if (reset) begin
      data_504 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_504 <= data_503;
        end
      end
    end
    if (reset) begin
      data_505 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_505 <= data_504;
        end
      end
    end
    if (reset) begin
      data_506 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_506 <= data_505;
        end
      end
    end
    if (reset) begin
      data_507 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_507 <= data_506;
        end
      end
    end
    if (reset) begin
      data_508 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_508 <= data_507;
        end
      end
    end
    if (reset) begin
      data_509 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_509 <= data_508;
        end
      end
    end
    if (reset) begin
      data_510 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_510 <= data_509;
        end
      end
    end
    if (reset) begin
      data_511 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_511 <= data_510;
        end
      end
    end
    if (reset) begin
      data_512 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_512 <= data_511;
        end
      end
    end
    if (reset) begin
      data_513 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_513 <= data_512;
        end
      end
    end
    if (reset) begin
      data_514 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_514 <= data_513;
        end
      end
    end
    if (reset) begin
      data_515 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_515 <= data_514;
        end
      end
    end
    if (reset) begin
      data_516 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_516 <= data_515;
        end
      end
    end
    if (reset) begin
      data_517 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_517 <= data_516;
        end
      end
    end
    if (reset) begin
      data_518 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_518 <= data_517;
        end
      end
    end
    if (reset) begin
      data_519 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_519 <= data_518;
        end
      end
    end
    if (reset) begin
      data_520 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_520 <= data_519;
        end
      end
    end
    if (reset) begin
      data_521 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_521 <= data_520;
        end
      end
    end
    if (reset) begin
      data_522 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_522 <= data_521;
        end
      end
    end
    if (reset) begin
      data_523 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_523 <= data_522;
        end
      end
    end
    if (reset) begin
      data_524 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_524 <= data_523;
        end
      end
    end
    if (reset) begin
      data_525 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_525 <= data_524;
        end
      end
    end
    if (reset) begin
      data_526 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_526 <= data_525;
        end
      end
    end
    if (reset) begin
      data_527 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_527 <= data_526;
        end
      end
    end
    if (reset) begin
      data_528 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_528 <= data_527;
        end
      end
    end
    if (reset) begin
      data_529 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_529 <= data_528;
        end
      end
    end
    if (reset) begin
      data_530 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_530 <= data_529;
        end
      end
    end
    if (reset) begin
      data_531 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_531 <= data_530;
        end
      end
    end
    if (reset) begin
      data_532 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_532 <= data_531;
        end
      end
    end
    if (reset) begin
      data_533 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_533 <= data_532;
        end
      end
    end
    if (reset) begin
      data_534 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_534 <= data_533;
        end
      end
    end
    if (reset) begin
      data_535 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_535 <= data_534;
        end
      end
    end
    if (reset) begin
      data_536 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_536 <= data_535;
        end
      end
    end
    if (reset) begin
      data_537 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_537 <= data_536;
        end
      end
    end
    if (reset) begin
      data_538 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_538 <= data_537;
        end
      end
    end
    if (reset) begin
      data_539 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_539 <= data_538;
        end
      end
    end
    if (reset) begin
      data_540 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_540 <= data_539;
        end
      end
    end
    if (reset) begin
      data_541 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_541 <= data_540;
        end
      end
    end
    if (reset) begin
      data_542 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_542 <= data_541;
        end
      end
    end
    if (reset) begin
      data_543 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_543 <= data_542;
        end
      end
    end
    if (reset) begin
      data_544 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_544 <= data_543;
        end
      end
    end
    if (reset) begin
      data_545 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_545 <= data_544;
        end
      end
    end
    if (reset) begin
      data_546 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_546 <= data_545;
        end
      end
    end
    if (reset) begin
      data_547 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_547 <= data_546;
        end
      end
    end
    if (reset) begin
      data_548 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_548 <= data_547;
        end
      end
    end
    if (reset) begin
      data_549 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_549 <= data_548;
        end
      end
    end
    if (reset) begin
      data_550 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_550 <= data_549;
        end
      end
    end
    if (reset) begin
      data_551 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_551 <= data_550;
        end
      end
    end
    if (reset) begin
      data_552 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_552 <= data_551;
        end
      end
    end
    if (reset) begin
      data_553 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_553 <= data_552;
        end
      end
    end
    if (reset) begin
      data_554 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_554 <= data_553;
        end
      end
    end
    if (reset) begin
      data_555 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_555 <= data_554;
        end
      end
    end
    if (reset) begin
      data_556 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_556 <= data_555;
        end
      end
    end
    if (reset) begin
      data_557 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_557 <= data_556;
        end
      end
    end
    if (reset) begin
      data_558 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_558 <= data_557;
        end
      end
    end
    if (reset) begin
      data_559 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_559 <= data_558;
        end
      end
    end
    if (reset) begin
      data_560 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_560 <= data_559;
        end
      end
    end
    if (reset) begin
      data_561 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_561 <= data_560;
        end
      end
    end
    if (reset) begin
      data_562 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_562 <= data_561;
        end
      end
    end
    if (reset) begin
      data_563 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_563 <= data_562;
        end
      end
    end
    if (reset) begin
      data_564 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_564 <= data_563;
        end
      end
    end
    if (reset) begin
      data_565 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_565 <= data_564;
        end
      end
    end
    if (reset) begin
      data_566 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_566 <= data_565;
        end
      end
    end
    if (reset) begin
      data_567 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_567 <= data_566;
        end
      end
    end
    if (reset) begin
      data_568 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_568 <= data_567;
        end
      end
    end
    if (reset) begin
      data_569 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_569 <= data_568;
        end
      end
    end
    if (reset) begin
      data_570 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_570 <= data_569;
        end
      end
    end
    if (reset) begin
      data_571 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_571 <= data_570;
        end
      end
    end
    if (reset) begin
      data_572 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_572 <= data_571;
        end
      end
    end
    if (reset) begin
      data_573 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_573 <= data_572;
        end
      end
    end
    if (reset) begin
      data_574 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_574 <= data_573;
        end
      end
    end
    if (reset) begin
      data_575 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_575 <= data_574;
        end
      end
    end
    if (reset) begin
      data_576 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_576 <= data_575;
        end
      end
    end
    if (reset) begin
      data_577 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_577 <= data_576;
        end
      end
    end
    if (reset) begin
      data_578 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_578 <= data_577;
        end
      end
    end
    if (reset) begin
      data_579 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_579 <= data_578;
        end
      end
    end
    if (reset) begin
      data_580 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_580 <= data_579;
        end
      end
    end
    if (reset) begin
      data_581 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_581 <= data_580;
        end
      end
    end
    if (reset) begin
      data_582 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_582 <= data_581;
        end
      end
    end
    if (reset) begin
      data_583 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_583 <= data_582;
        end
      end
    end
    if (reset) begin
      data_584 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_584 <= data_583;
        end
      end
    end
    if (reset) begin
      data_585 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_585 <= data_584;
        end
      end
    end
    if (reset) begin
      data_586 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_586 <= data_585;
        end
      end
    end
    if (reset) begin
      data_587 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_587 <= data_586;
        end
      end
    end
    if (reset) begin
      data_588 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_588 <= data_587;
        end
      end
    end
    if (reset) begin
      data_589 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_589 <= data_588;
        end
      end
    end
    if (reset) begin
      data_590 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_590 <= data_589;
        end
      end
    end
    if (reset) begin
      data_591 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_591 <= data_590;
        end
      end
    end
    if (reset) begin
      data_592 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_592 <= data_591;
        end
      end
    end
    if (reset) begin
      data_593 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_593 <= data_592;
        end
      end
    end
    if (reset) begin
      data_594 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_594 <= data_593;
        end
      end
    end
    if (reset) begin
      data_595 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_595 <= data_594;
        end
      end
    end
    if (reset) begin
      data_596 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_596 <= data_595;
        end
      end
    end
    if (reset) begin
      data_597 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_597 <= data_596;
        end
      end
    end
    if (reset) begin
      data_598 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_598 <= data_597;
        end
      end
    end
    if (reset) begin
      data_599 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_599 <= data_598;
        end
      end
    end
    if (reset) begin
      data_600 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_600 <= data_599;
        end
      end
    end
    if (reset) begin
      data_601 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_601 <= data_600;
        end
      end
    end
    if (reset) begin
      data_602 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_602 <= data_601;
        end
      end
    end
    if (reset) begin
      data_603 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_603 <= data_602;
        end
      end
    end
    if (reset) begin
      data_604 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_604 <= data_603;
        end
      end
    end
    if (reset) begin
      data_605 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_605 <= data_604;
        end
      end
    end
    if (reset) begin
      data_606 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_606 <= data_605;
        end
      end
    end
    if (reset) begin
      data_607 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_607 <= data_606;
        end
      end
    end
    if (reset) begin
      data_608 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_608 <= data_607;
        end
      end
    end
    if (reset) begin
      data_609 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_609 <= data_608;
        end
      end
    end
    if (reset) begin
      data_610 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_610 <= data_609;
        end
      end
    end
    if (reset) begin
      data_611 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_611 <= data_610;
        end
      end
    end
    if (reset) begin
      data_612 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_612 <= data_611;
        end
      end
    end
    if (reset) begin
      data_613 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_613 <= data_612;
        end
      end
    end
    if (reset) begin
      data_614 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_614 <= data_613;
        end
      end
    end
    if (reset) begin
      data_615 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_615 <= data_614;
        end
      end
    end
    if (reset) begin
      data_616 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_616 <= data_615;
        end
      end
    end
    if (reset) begin
      data_617 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_617 <= data_616;
        end
      end
    end
    if (reset) begin
      data_618 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_618 <= data_617;
        end
      end
    end
    if (reset) begin
      data_619 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_619 <= data_618;
        end
      end
    end
    if (reset) begin
      data_620 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_620 <= data_619;
        end
      end
    end
    if (reset) begin
      data_621 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_621 <= data_620;
        end
      end
    end
    if (reset) begin
      data_622 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_622 <= data_621;
        end
      end
    end
    if (reset) begin
      data_623 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_623 <= data_622;
        end
      end
    end
    if (reset) begin
      data_624 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_624 <= data_623;
        end
      end
    end
    if (reset) begin
      data_625 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_625 <= data_624;
        end
      end
    end
    if (reset) begin
      data_626 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_626 <= data_625;
        end
      end
    end
    if (reset) begin
      data_627 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_627 <= data_626;
        end
      end
    end
    if (reset) begin
      data_628 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_628 <= data_627;
        end
      end
    end
    if (reset) begin
      data_629 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_629 <= data_628;
        end
      end
    end
    if (reset) begin
      data_630 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_630 <= data_629;
        end
      end
    end
    if (reset) begin
      data_631 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_631 <= data_630;
        end
      end
    end
    if (reset) begin
      data_632 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_632 <= data_631;
        end
      end
    end
    if (reset) begin
      data_633 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_633 <= data_632;
        end
      end
    end
    if (reset) begin
      data_634 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_634 <= data_633;
        end
      end
    end
    if (reset) begin
      data_635 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_635 <= data_634;
        end
      end
    end
    if (reset) begin
      data_636 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_636 <= data_635;
        end
      end
    end
    if (reset) begin
      data_637 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_637 <= data_636;
        end
      end
    end
    if (reset) begin
      data_638 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_638 <= data_637;
        end
      end
    end
    if (reset) begin
      data_639 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_639 <= data_638;
        end
      end
    end
    if (reset) begin
      data_640 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_640 <= data_639;
        end
      end
    end
    if (reset) begin
      data_641 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_641 <= data_640;
        end
      end
    end
    if (reset) begin
      data_642 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_642 <= data_641;
        end
      end
    end
    if (reset) begin
      data_643 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_643 <= data_642;
        end
      end
    end
    if (reset) begin
      data_644 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_644 <= data_643;
        end
      end
    end
    if (reset) begin
      data_645 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_645 <= data_644;
        end
      end
    end
    if (reset) begin
      data_646 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_646 <= data_645;
        end
      end
    end
    if (reset) begin
      data_647 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_647 <= data_646;
        end
      end
    end
    if (reset) begin
      data_648 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_648 <= data_647;
        end
      end
    end
    if (reset) begin
      data_649 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_649 <= data_648;
        end
      end
    end
    if (reset) begin
      data_650 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_650 <= data_649;
        end
      end
    end
    if (reset) begin
      data_651 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_651 <= data_650;
        end
      end
    end
    if (reset) begin
      data_652 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_652 <= data_651;
        end
      end
    end
    if (reset) begin
      data_653 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_653 <= data_652;
        end
      end
    end
    if (reset) begin
      data_654 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_654 <= data_653;
        end
      end
    end
    if (reset) begin
      data_655 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_655 <= data_654;
        end
      end
    end
    if (reset) begin
      data_656 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_656 <= data_655;
        end
      end
    end
    if (reset) begin
      data_657 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_657 <= data_656;
        end
      end
    end
    if (reset) begin
      data_658 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_658 <= data_657;
        end
      end
    end
    if (reset) begin
      data_659 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_659 <= data_658;
        end
      end
    end
    if (reset) begin
      data_660 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_660 <= data_659;
        end
      end
    end
    if (reset) begin
      data_661 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_661 <= data_660;
        end
      end
    end
    if (reset) begin
      data_662 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_662 <= data_661;
        end
      end
    end
    if (reset) begin
      data_663 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_663 <= data_662;
        end
      end
    end
    if (reset) begin
      data_664 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_664 <= data_663;
        end
      end
    end
    if (reset) begin
      data_665 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_665 <= data_664;
        end
      end
    end
    if (reset) begin
      data_666 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_666 <= data_665;
        end
      end
    end
    if (reset) begin
      data_667 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_667 <= data_666;
        end
      end
    end
    if (reset) begin
      data_668 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_668 <= data_667;
        end
      end
    end
    if (reset) begin
      data_669 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_669 <= data_668;
        end
      end
    end
    if (reset) begin
      data_670 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_670 <= data_669;
        end
      end
    end
    if (reset) begin
      data_671 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_671 <= data_670;
        end
      end
    end
    if (reset) begin
      data_672 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_672 <= data_671;
        end
      end
    end
    if (reset) begin
      data_673 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_673 <= data_672;
        end
      end
    end
    if (reset) begin
      data_674 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_674 <= data_673;
        end
      end
    end
    if (reset) begin
      data_675 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_675 <= data_674;
        end
      end
    end
    if (reset) begin
      data_676 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_676 <= data_675;
        end
      end
    end
    if (reset) begin
      data_677 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_677 <= data_676;
        end
      end
    end
    if (reset) begin
      data_678 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_678 <= data_677;
        end
      end
    end
    if (reset) begin
      data_679 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_679 <= data_678;
        end
      end
    end
    if (reset) begin
      data_680 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_680 <= data_679;
        end
      end
    end
    if (reset) begin
      data_681 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_681 <= data_680;
        end
      end
    end
    if (reset) begin
      data_682 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_682 <= data_681;
        end
      end
    end
    if (reset) begin
      data_683 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_683 <= data_682;
        end
      end
    end
    if (reset) begin
      data_684 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_684 <= data_683;
        end
      end
    end
    if (reset) begin
      data_685 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_685 <= data_684;
        end
      end
    end
    if (reset) begin
      data_686 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_686 <= data_685;
        end
      end
    end
    if (reset) begin
      data_687 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_687 <= data_686;
        end
      end
    end
    if (reset) begin
      data_688 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_688 <= data_687;
        end
      end
    end
    if (reset) begin
      data_689 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_689 <= data_688;
        end
      end
    end
    if (reset) begin
      data_690 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_690 <= data_689;
        end
      end
    end
    if (reset) begin
      data_691 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_691 <= data_690;
        end
      end
    end
    if (reset) begin
      data_692 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_692 <= data_691;
        end
      end
    end
    if (reset) begin
      data_693 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_693 <= data_692;
        end
      end
    end
    if (reset) begin
      data_694 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_694 <= data_693;
        end
      end
    end
    if (reset) begin
      data_695 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_695 <= data_694;
        end
      end
    end
    if (reset) begin
      data_696 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_696 <= data_695;
        end
      end
    end
    if (reset) begin
      data_697 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_697 <= data_696;
        end
      end
    end
    if (reset) begin
      data_698 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_698 <= data_697;
        end
      end
    end
    if (reset) begin
      data_699 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_699 <= data_698;
        end
      end
    end
    if (reset) begin
      data_700 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_700 <= data_699;
        end
      end
    end
    if (reset) begin
      data_701 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_701 <= data_700;
        end
      end
    end
    if (reset) begin
      data_702 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_702 <= data_701;
        end
      end
    end
    if (reset) begin
      data_703 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_703 <= data_702;
        end
      end
    end
    if (reset) begin
      data_704 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_704 <= data_703;
        end
      end
    end
    if (reset) begin
      data_705 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_705 <= data_704;
        end
      end
    end
    if (reset) begin
      data_706 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_706 <= data_705;
        end
      end
    end
    if (reset) begin
      data_707 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_707 <= data_706;
        end
      end
    end
    if (reset) begin
      data_708 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_708 <= data_707;
        end
      end
    end
    if (reset) begin
      data_709 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_709 <= data_708;
        end
      end
    end
    if (reset) begin
      data_710 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_710 <= data_709;
        end
      end
    end
    if (reset) begin
      data_711 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_711 <= data_710;
        end
      end
    end
    if (reset) begin
      data_712 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_712 <= data_711;
        end
      end
    end
    if (reset) begin
      data_713 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_713 <= data_712;
        end
      end
    end
    if (reset) begin
      data_714 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_714 <= data_713;
        end
      end
    end
    if (reset) begin
      data_715 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_715 <= data_714;
        end
      end
    end
    if (reset) begin
      data_716 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_716 <= data_715;
        end
      end
    end
    if (reset) begin
      data_717 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_717 <= data_716;
        end
      end
    end
    if (reset) begin
      data_718 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_718 <= data_717;
        end
      end
    end
    if (reset) begin
      data_719 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_719 <= data_718;
        end
      end
    end
    if (reset) begin
      data_720 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_720 <= data_719;
        end
      end
    end
    if (reset) begin
      data_721 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_721 <= data_720;
        end
      end
    end
    if (reset) begin
      data_722 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_722 <= data_721;
        end
      end
    end
    if (reset) begin
      data_723 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_723 <= data_722;
        end
      end
    end
    if (reset) begin
      data_724 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_724 <= data_723;
        end
      end
    end
    if (reset) begin
      data_725 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_725 <= data_724;
        end
      end
    end
    if (reset) begin
      data_726 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_726 <= data_725;
        end
      end
    end
    if (reset) begin
      data_727 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_727 <= data_726;
        end
      end
    end
    if (reset) begin
      data_728 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_728 <= data_727;
        end
      end
    end
    if (reset) begin
      data_729 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_729 <= data_728;
        end
      end
    end
    if (reset) begin
      data_730 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_730 <= data_729;
        end
      end
    end
    if (reset) begin
      data_731 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_731 <= data_730;
        end
      end
    end
    if (reset) begin
      data_732 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_732 <= data_731;
        end
      end
    end
    if (reset) begin
      data_733 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_733 <= data_732;
        end
      end
    end
    if (reset) begin
      data_734 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_734 <= data_733;
        end
      end
    end
    if (reset) begin
      data_735 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_735 <= data_734;
        end
      end
    end
    if (reset) begin
      data_736 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_736 <= data_735;
        end
      end
    end
    if (reset) begin
      data_737 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_737 <= data_736;
        end
      end
    end
    if (reset) begin
      data_738 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_738 <= data_737;
        end
      end
    end
    if (reset) begin
      data_739 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_739 <= data_738;
        end
      end
    end
    if (reset) begin
      data_740 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_740 <= data_739;
        end
      end
    end
    if (reset) begin
      data_741 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_741 <= data_740;
        end
      end
    end
    if (reset) begin
      data_742 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_742 <= data_741;
        end
      end
    end
    if (reset) begin
      data_743 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_743 <= data_742;
        end
      end
    end
    if (reset) begin
      data_744 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_744 <= data_743;
        end
      end
    end
    if (reset) begin
      data_745 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_745 <= data_744;
        end
      end
    end
    if (reset) begin
      data_746 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_746 <= data_745;
        end
      end
    end
    if (reset) begin
      data_747 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_747 <= data_746;
        end
      end
    end
    if (reset) begin
      data_748 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_748 <= data_747;
        end
      end
    end
    if (reset) begin
      data_749 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_749 <= data_748;
        end
      end
    end
    if (reset) begin
      data_750 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_750 <= data_749;
        end
      end
    end
    if (reset) begin
      data_751 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_751 <= data_750;
        end
      end
    end
    if (reset) begin
      data_752 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_752 <= data_751;
        end
      end
    end
    if (reset) begin
      data_753 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_753 <= data_752;
        end
      end
    end
    if (reset) begin
      data_754 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_754 <= data_753;
        end
      end
    end
    if (reset) begin
      data_755 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_755 <= data_754;
        end
      end
    end
    if (reset) begin
      data_756 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_756 <= data_755;
        end
      end
    end
    if (reset) begin
      data_757 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_757 <= data_756;
        end
      end
    end
    if (reset) begin
      data_758 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_758 <= data_757;
        end
      end
    end
    if (reset) begin
      data_759 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_759 <= data_758;
        end
      end
    end
    if (reset) begin
      data_760 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_760 <= data_759;
        end
      end
    end
    if (reset) begin
      data_761 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_761 <= data_760;
        end
      end
    end
    if (reset) begin
      data_762 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_762 <= data_761;
        end
      end
    end
    if (reset) begin
      data_763 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_763 <= data_762;
        end
      end
    end
    if (reset) begin
      data_764 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_764 <= data_763;
        end
      end
    end
    if (reset) begin
      data_765 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_765 <= data_764;
        end
      end
    end
    if (reset) begin
      data_766 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_766 <= data_765;
        end
      end
    end
    if (reset) begin
      data_767 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_767 <= data_766;
        end
      end
    end
    if (reset) begin
      data_768 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_768 <= data_767;
        end
      end
    end
    if (reset) begin
      data_769 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_769 <= data_768;
        end
      end
    end
    if (reset) begin
      data_770 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_770 <= data_769;
        end
      end
    end
    if (reset) begin
      data_771 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_771 <= data_770;
        end
      end
    end
    if (reset) begin
      data_772 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_772 <= data_771;
        end
      end
    end
    if (reset) begin
      data_773 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_773 <= data_772;
        end
      end
    end
    if (reset) begin
      data_774 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_774 <= data_773;
        end
      end
    end
    if (reset) begin
      data_775 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_775 <= data_774;
        end
      end
    end
    if (reset) begin
      data_776 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_776 <= data_775;
        end
      end
    end
    if (reset) begin
      data_777 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_777 <= data_776;
        end
      end
    end
    if (reset) begin
      data_778 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_778 <= data_777;
        end
      end
    end
    if (reset) begin
      data_779 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_779 <= data_778;
        end
      end
    end
    if (reset) begin
      data_780 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_780 <= data_779;
        end
      end
    end
    if (reset) begin
      data_781 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_781 <= data_780;
        end
      end
    end
    if (reset) begin
      data_782 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_782 <= data_781;
        end
      end
    end
    if (reset) begin
      data_783 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_783 <= data_782;
        end
      end
    end
    if (reset) begin
      data_784 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_784 <= data_783;
        end
      end
    end
    if (reset) begin
      data_785 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_785 <= data_784;
        end
      end
    end
    if (reset) begin
      data_786 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_786 <= data_785;
        end
      end
    end
    if (reset) begin
      data_787 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_787 <= data_786;
        end
      end
    end
    if (reset) begin
      data_788 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_788 <= data_787;
        end
      end
    end
    if (reset) begin
      data_789 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_789 <= data_788;
        end
      end
    end
    if (reset) begin
      data_790 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_790 <= data_789;
        end
      end
    end
    if (reset) begin
      data_791 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_791 <= data_790;
        end
      end
    end
    if (reset) begin
      data_792 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_792 <= data_791;
        end
      end
    end
    if (reset) begin
      data_793 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_793 <= data_792;
        end
      end
    end
    if (reset) begin
      data_794 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_794 <= data_793;
        end
      end
    end
    if (reset) begin
      data_795 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_795 <= data_794;
        end
      end
    end
    if (reset) begin
      data_796 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_796 <= data_795;
        end
      end
    end
    if (reset) begin
      data_797 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_797 <= data_796;
        end
      end
    end
    if (reset) begin
      data_798 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_798 <= data_797;
        end
      end
    end
    if (reset) begin
      data_799 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_799 <= data_798;
        end
      end
    end
    if (reset) begin
      data_800 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_800 <= data_799;
        end
      end
    end
    if (reset) begin
      data_801 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_801 <= data_800;
        end
      end
    end
    if (reset) begin
      data_802 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_802 <= data_801;
        end
      end
    end
    if (reset) begin
      data_803 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_803 <= data_802;
        end
      end
    end
    if (reset) begin
      data_804 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_804 <= data_803;
        end
      end
    end
    if (reset) begin
      data_805 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_805 <= data_804;
        end
      end
    end
    if (reset) begin
      data_806 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_806 <= data_805;
        end
      end
    end
    if (reset) begin
      data_807 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_807 <= data_806;
        end
      end
    end
    if (reset) begin
      data_808 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_808 <= data_807;
        end
      end
    end
    if (reset) begin
      data_809 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_809 <= data_808;
        end
      end
    end
    if (reset) begin
      data_810 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_810 <= data_809;
        end
      end
    end
    if (reset) begin
      data_811 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_811 <= data_810;
        end
      end
    end
    if (reset) begin
      data_812 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_812 <= data_811;
        end
      end
    end
    if (reset) begin
      data_813 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_813 <= data_812;
        end
      end
    end
    if (reset) begin
      data_814 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_814 <= data_813;
        end
      end
    end
    if (reset) begin
      data_815 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_815 <= data_814;
        end
      end
    end
    if (reset) begin
      data_816 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_816 <= data_815;
        end
      end
    end
    if (reset) begin
      data_817 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_817 <= data_816;
        end
      end
    end
    if (reset) begin
      data_818 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_818 <= data_817;
        end
      end
    end
    if (reset) begin
      data_819 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_819 <= data_818;
        end
      end
    end
    if (reset) begin
      data_820 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_820 <= data_819;
        end
      end
    end
    if (reset) begin
      data_821 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_821 <= data_820;
        end
      end
    end
    if (reset) begin
      data_822 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_822 <= data_821;
        end
      end
    end
    if (reset) begin
      data_823 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_823 <= data_822;
        end
      end
    end
    if (reset) begin
      data_824 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_824 <= data_823;
        end
      end
    end
    if (reset) begin
      data_825 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_825 <= data_824;
        end
      end
    end
    if (reset) begin
      data_826 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_826 <= data_825;
        end
      end
    end
    if (reset) begin
      data_827 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_827 <= data_826;
        end
      end
    end
    if (reset) begin
      data_828 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_828 <= data_827;
        end
      end
    end
    if (reset) begin
      data_829 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_829 <= data_828;
        end
      end
    end
    if (reset) begin
      data_830 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_830 <= data_829;
        end
      end
    end
    if (reset) begin
      data_831 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_831 <= data_830;
        end
      end
    end
    if (reset) begin
      data_832 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_832 <= data_831;
        end
      end
    end
    if (reset) begin
      data_833 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_833 <= data_832;
        end
      end
    end
    if (reset) begin
      data_834 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_834 <= data_833;
        end
      end
    end
    if (reset) begin
      data_835 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_835 <= data_834;
        end
      end
    end
    if (reset) begin
      data_836 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_836 <= data_835;
        end
      end
    end
    if (reset) begin
      data_837 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_837 <= data_836;
        end
      end
    end
    if (reset) begin
      data_838 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_838 <= data_837;
        end
      end
    end
    if (reset) begin
      data_839 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_839 <= data_838;
        end
      end
    end
    if (reset) begin
      data_840 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_840 <= data_839;
        end
      end
    end
    if (reset) begin
      data_841 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_841 <= data_840;
        end
      end
    end
    if (reset) begin
      data_842 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_842 <= data_841;
        end
      end
    end
    if (reset) begin
      data_843 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_843 <= data_842;
        end
      end
    end
    if (reset) begin
      data_844 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_844 <= data_843;
        end
      end
    end
    if (reset) begin
      data_845 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_845 <= data_844;
        end
      end
    end
    if (reset) begin
      data_846 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_846 <= data_845;
        end
      end
    end
    if (reset) begin
      data_847 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_847 <= data_846;
        end
      end
    end
    if (reset) begin
      data_848 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_848 <= data_847;
        end
      end
    end
    if (reset) begin
      data_849 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_849 <= data_848;
        end
      end
    end
    if (reset) begin
      data_850 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_850 <= data_849;
        end
      end
    end
    if (reset) begin
      data_851 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_851 <= data_850;
        end
      end
    end
    if (reset) begin
      data_852 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_852 <= data_851;
        end
      end
    end
    if (reset) begin
      data_853 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_853 <= data_852;
        end
      end
    end
    if (reset) begin
      data_854 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_854 <= data_853;
        end
      end
    end
    if (reset) begin
      data_855 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_855 <= data_854;
        end
      end
    end
    if (reset) begin
      data_856 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_856 <= data_855;
        end
      end
    end
    if (reset) begin
      data_857 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_857 <= data_856;
        end
      end
    end
    if (reset) begin
      data_858 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_858 <= data_857;
        end
      end
    end
    if (reset) begin
      data_859 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_859 <= data_858;
        end
      end
    end
    if (reset) begin
      data_860 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_860 <= data_859;
        end
      end
    end
    if (reset) begin
      data_861 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_861 <= data_860;
        end
      end
    end
    if (reset) begin
      data_862 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_862 <= data_861;
        end
      end
    end
    if (reset) begin
      data_863 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_863 <= data_862;
        end
      end
    end
    if (reset) begin
      data_864 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_864 <= data_863;
        end
      end
    end
    if (reset) begin
      data_865 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_865 <= data_864;
        end
      end
    end
    if (reset) begin
      data_866 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_866 <= data_865;
        end
      end
    end
    if (reset) begin
      data_867 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_867 <= data_866;
        end
      end
    end
    if (reset) begin
      data_868 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_868 <= data_867;
        end
      end
    end
    if (reset) begin
      data_869 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_869 <= data_868;
        end
      end
    end
    if (reset) begin
      data_870 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_870 <= data_869;
        end
      end
    end
    if (reset) begin
      data_871 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_871 <= data_870;
        end
      end
    end
    if (reset) begin
      data_872 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_872 <= data_871;
        end
      end
    end
    if (reset) begin
      data_873 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_873 <= data_872;
        end
      end
    end
    if (reset) begin
      data_874 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_874 <= data_873;
        end
      end
    end
    if (reset) begin
      data_875 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_875 <= data_874;
        end
      end
    end
    if (reset) begin
      data_876 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_876 <= data_875;
        end
      end
    end
    if (reset) begin
      data_877 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_877 <= data_876;
        end
      end
    end
    if (reset) begin
      data_878 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_878 <= data_877;
        end
      end
    end
    if (reset) begin
      data_879 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_879 <= data_878;
        end
      end
    end
    if (reset) begin
      data_880 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_880 <= data_879;
        end
      end
    end
    if (reset) begin
      data_881 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_881 <= data_880;
        end
      end
    end
    if (reset) begin
      data_882 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_882 <= data_881;
        end
      end
    end
    if (reset) begin
      data_883 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_883 <= data_882;
        end
      end
    end
    if (reset) begin
      data_884 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_884 <= data_883;
        end
      end
    end
    if (reset) begin
      data_885 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_885 <= data_884;
        end
      end
    end
    if (reset) begin
      data_886 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_886 <= data_885;
        end
      end
    end
    if (reset) begin
      data_887 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_887 <= data_886;
        end
      end
    end
    if (reset) begin
      data_888 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_888 <= data_887;
        end
      end
    end
    if (reset) begin
      data_889 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_889 <= data_888;
        end
      end
    end
    if (reset) begin
      data_890 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_890 <= data_889;
        end
      end
    end
    if (reset) begin
      data_891 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_891 <= data_890;
        end
      end
    end
    if (reset) begin
      data_892 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_892 <= data_891;
        end
      end
    end
    if (reset) begin
      data_893 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_893 <= data_892;
        end
      end
    end
    if (reset) begin
      data_894 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_894 <= data_893;
        end
      end
    end
    if (reset) begin
      data_895 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_895 <= data_894;
        end
      end
    end
    if (reset) begin
      data_896 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_896 <= data_895;
        end
      end
    end
    if (reset) begin
      data_897 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_897 <= data_896;
        end
      end
    end
    if (reset) begin
      data_898 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_898 <= data_897;
        end
      end
    end
    if (reset) begin
      data_899 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_899 <= data_898;
        end
      end
    end
    if (reset) begin
      data_900 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_900 <= data_899;
        end
      end
    end
    if (reset) begin
      data_901 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_901 <= data_900;
        end
      end
    end
    if (reset) begin
      data_902 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_902 <= data_901;
        end
      end
    end
    if (reset) begin
      data_903 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_903 <= data_902;
        end
      end
    end
    if (reset) begin
      data_904 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_904 <= data_903;
        end
      end
    end
    if (reset) begin
      data_905 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_905 <= data_904;
        end
      end
    end
    if (reset) begin
      data_906 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_906 <= data_905;
        end
      end
    end
    if (reset) begin
      data_907 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_907 <= data_906;
        end
      end
    end
    if (reset) begin
      data_908 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_908 <= data_907;
        end
      end
    end
    if (reset) begin
      data_909 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_909 <= data_908;
        end
      end
    end
    if (reset) begin
      data_910 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_910 <= data_909;
        end
      end
    end
    if (reset) begin
      data_911 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_911 <= data_910;
        end
      end
    end
    if (reset) begin
      data_912 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_912 <= data_911;
        end
      end
    end
    if (reset) begin
      data_913 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_913 <= data_912;
        end
      end
    end
    if (reset) begin
      data_914 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_914 <= data_913;
        end
      end
    end
    if (reset) begin
      data_915 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_915 <= data_914;
        end
      end
    end
    if (reset) begin
      data_916 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_916 <= data_915;
        end
      end
    end
    if (reset) begin
      data_917 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_917 <= data_916;
        end
      end
    end
    if (reset) begin
      data_918 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_918 <= data_917;
        end
      end
    end
    if (reset) begin
      data_919 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_919 <= data_918;
        end
      end
    end
    if (reset) begin
      data_920 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_920 <= data_919;
        end
      end
    end
    if (reset) begin
      data_921 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_921 <= data_920;
        end
      end
    end
    if (reset) begin
      data_922 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_922 <= data_921;
        end
      end
    end
    if (reset) begin
      data_923 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_923 <= data_922;
        end
      end
    end
    if (reset) begin
      data_924 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_924 <= data_923;
        end
      end
    end
    if (reset) begin
      data_925 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_925 <= data_924;
        end
      end
    end
    if (reset) begin
      data_926 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_926 <= data_925;
        end
      end
    end
    if (reset) begin
      data_927 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_927 <= data_926;
        end
      end
    end
    if (reset) begin
      data_928 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_928 <= data_927;
        end
      end
    end
    if (reset) begin
      data_929 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_929 <= data_928;
        end
      end
    end
    if (reset) begin
      data_930 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_930 <= data_929;
        end
      end
    end
    if (reset) begin
      data_931 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_931 <= data_930;
        end
      end
    end
    if (reset) begin
      data_932 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_932 <= data_931;
        end
      end
    end
    if (reset) begin
      data_933 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_933 <= data_932;
        end
      end
    end
    if (reset) begin
      data_934 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_934 <= data_933;
        end
      end
    end
    if (reset) begin
      data_935 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_935 <= data_934;
        end
      end
    end
    if (reset) begin
      data_936 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_936 <= data_935;
        end
      end
    end
    if (reset) begin
      data_937 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_937 <= data_936;
        end
      end
    end
    if (reset) begin
      data_938 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_938 <= data_937;
        end
      end
    end
    if (reset) begin
      data_939 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_939 <= data_938;
        end
      end
    end
    if (reset) begin
      data_940 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_940 <= data_939;
        end
      end
    end
    if (reset) begin
      data_941 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_941 <= data_940;
        end
      end
    end
    if (reset) begin
      data_942 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_942 <= data_941;
        end
      end
    end
    if (reset) begin
      data_943 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_943 <= data_942;
        end
      end
    end
    if (reset) begin
      data_944 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_944 <= data_943;
        end
      end
    end
    if (reset) begin
      data_945 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_945 <= data_944;
        end
      end
    end
    if (reset) begin
      data_946 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_946 <= data_945;
        end
      end
    end
    if (reset) begin
      data_947 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_947 <= data_946;
        end
      end
    end
    if (reset) begin
      data_948 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_948 <= data_947;
        end
      end
    end
    if (reset) begin
      data_949 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_949 <= data_948;
        end
      end
    end
    if (reset) begin
      data_950 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_950 <= data_949;
        end
      end
    end
    if (reset) begin
      data_951 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_951 <= data_950;
        end
      end
    end
    if (reset) begin
      data_952 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_952 <= data_951;
        end
      end
    end
    if (reset) begin
      data_953 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_953 <= data_952;
        end
      end
    end
    if (reset) begin
      data_954 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_954 <= data_953;
        end
      end
    end
    if (reset) begin
      data_955 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_955 <= data_954;
        end
      end
    end
    if (reset) begin
      data_956 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_956 <= data_955;
        end
      end
    end
    if (reset) begin
      data_957 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_957 <= data_956;
        end
      end
    end
    if (reset) begin
      data_958 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_958 <= data_957;
        end
      end
    end
    if (reset) begin
      data_959 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_959 <= data_958;
        end
      end
    end
    if (reset) begin
      data_960 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_960 <= data_959;
        end
      end
    end
    if (reset) begin
      data_961 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_961 <= data_960;
        end
      end
    end
    if (reset) begin
      data_962 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_962 <= data_961;
        end
      end
    end
    if (reset) begin
      data_963 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_963 <= data_962;
        end
      end
    end
    if (reset) begin
      data_964 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_964 <= data_963;
        end
      end
    end
    if (reset) begin
      data_965 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_965 <= data_964;
        end
      end
    end
    if (reset) begin
      data_966 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_966 <= data_965;
        end
      end
    end
    if (reset) begin
      data_967 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_967 <= data_966;
        end
      end
    end
    if (reset) begin
      data_968 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_968 <= data_967;
        end
      end
    end
    if (reset) begin
      data_969 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_969 <= data_968;
        end
      end
    end
    if (reset) begin
      data_970 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_970 <= data_969;
        end
      end
    end
    if (reset) begin
      data_971 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_971 <= data_970;
        end
      end
    end
    if (reset) begin
      data_972 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_972 <= data_971;
        end
      end
    end
    if (reset) begin
      data_973 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_973 <= data_972;
        end
      end
    end
    if (reset) begin
      data_974 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_974 <= data_973;
        end
      end
    end
    if (reset) begin
      data_975 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_975 <= data_974;
        end
      end
    end
    if (reset) begin
      data_976 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_976 <= data_975;
        end
      end
    end
    if (reset) begin
      data_977 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_977 <= data_976;
        end
      end
    end
    if (reset) begin
      data_978 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_978 <= data_977;
        end
      end
    end
    if (reset) begin
      data_979 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_979 <= data_978;
        end
      end
    end
    if (reset) begin
      data_980 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_980 <= data_979;
        end
      end
    end
    if (reset) begin
      data_981 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_981 <= data_980;
        end
      end
    end
    if (reset) begin
      data_982 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_982 <= data_981;
        end
      end
    end
    if (reset) begin
      data_983 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_983 <= data_982;
        end
      end
    end
    if (reset) begin
      data_984 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_984 <= data_983;
        end
      end
    end
    if (reset) begin
      data_985 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_985 <= data_984;
        end
      end
    end
    if (reset) begin
      data_986 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_986 <= data_985;
        end
      end
    end
    if (reset) begin
      data_987 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_987 <= data_986;
        end
      end
    end
    if (reset) begin
      data_988 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_988 <= data_987;
        end
      end
    end
    if (reset) begin
      data_989 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_989 <= data_988;
        end
      end
    end
    if (reset) begin
      data_990 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_990 <= data_989;
        end
      end
    end
    if (reset) begin
      data_991 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_991 <= data_990;
        end
      end
    end
    if (reset) begin
      data_992 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_992 <= data_991;
        end
      end
    end
    if (reset) begin
      data_993 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_993 <= data_992;
        end
      end
    end
    if (reset) begin
      data_994 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_994 <= data_993;
        end
      end
    end
    if (reset) begin
      data_995 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_995 <= data_994;
        end
      end
    end
    if (reset) begin
      data_996 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_996 <= data_995;
        end
      end
    end
    if (reset) begin
      data_997 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_997 <= data_996;
        end
      end
    end
    if (reset) begin
      data_998 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_998 <= data_997;
        end
      end
    end
    if (reset) begin
      data_999 <= 32'sh0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_999 <= data_998;
        end
      end
    end
    if (reset) begin
      result <= 64'sh0;
    end else begin
      result <= _GEN_6003[79:16];
    end
  end
endmodule
