// SPDX-License-Identifier: Apache-2.0
// Example VCS Command: $VCS_HOME/bin/vcs -debug_pp -full64 +define+UNIT_DELAY +rad +v2k +vcs+lic+wait +vc+list +vcs+initreg+random +vcs+dumpvars+out.vcd tb.v SCIEPipelined.v ...
`timescale 100ps / 10ps

`define CLK_PERIOD 1

`define HALF_CLK_PERIOD 0.5
`define RESET_TIME 5
`define INIT_TIME 5.5
`define expect(nodeName, nodeVal, expVal, cycle) if (nodeVal !== expVal) begin \
  $display("\t ASSERTION ON %s FAILED @ CYCLE = %d, 0x%h != EXPECTED 0x%h", \
  nodeName,cycle,nodeVal,expVal); $stop; end

module testbench_v;

  integer cycle = 0;

  reg clock = 1;
  reg reset = 1;
  reg[31:0] io_rs2 = 0;
  reg signed [31:0] io_rs1 = 0;
  reg[31:0] io_insn = 0;
  reg[0:0] io_valid = 0;
  wire signed [31:0] io_rd;

  always #`HALF_CLK_PERIOD clock = ~clock;

  initial begin
    #`RESET_TIME
    forever #`CLK_PERIOD cycle = cycle + 1;
  end

  SCIEPipelined SCIEPipelined(
    .clock(clock),
    .reset(reset),
    .io_rs2(io_rs2),
    .io_rs1(io_rs1),
    .io_insn(io_insn),
    .io_valid(io_valid),
    .io_rd(io_rd));

  initial begin
    #`INIT_TIME reset = 0;
    io_valid = 1'd1;
    io_insn = 4'd11;
    io_rs1 = 22'd2727536;
    io_rs2 = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 4'd11;
    io_rs1 = 21'd1107598;
    io_rs2 = 1'd1;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 4'd11;
    io_rs1 = 23'd5162021;
    io_rs2 = 2'd2;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 4'd11;
    io_rs1 = 22'd2528178;
    io_rs2 = 2'd3;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 4'd11;
    io_rs1 = 22'd2760774;
    io_rs2 = 3'd4;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd6156421;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,256223448,cycle)
    `expect("io_rd",io_rd,256223448,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3047181;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,230867545,cycle)
    `expect("io_rd",io_rd,230867545,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 20'd838509;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,571314843,cycle)
    `expect("io_rd",io_rd,571314843,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 16'd42700;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,493459123,cycle)
    `expect("io_rd",io_rd,493459123,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2313773;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,539961206,cycle)
    `expect("io_rd",io_rd,539961206,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd4031849;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,370981445,cycle)
    `expect("io_rd",io_rd,370981445,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3646793;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,439133589,cycle)
    `expect("io_rd",io_rd,439133589,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 18'd168310;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,477268317,cycle)
    `expect("io_rd",io_rd,477268317,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 16'd43739;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,544915433,cycle)
    `expect("io_rd",io_rd,544915433,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 20'd964250;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,364655415,cycle)
    `expect("io_rd",io_rd,364655415,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5109807;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,392524024,cycle)
    `expect("io_rd",io_rd,392524024,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 19'd442457;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,189501251,cycle)
    `expect("io_rd",io_rd,189501251,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd4138661;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,621244682,cycle)
    `expect("io_rd",io_rd,621244682,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 20'd658333;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,369936369,cycle)
    `expect("io_rd",io_rd,369936369,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5349771;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,792089060,cycle)
    `expect("io_rd",io_rd,792089060,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5650834;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,555746049,cycle)
    `expect("io_rd",io_rd,555746049,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd6280114;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,977996984,cycle)
    `expect("io_rd",io_rd,977996984,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3388914;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,926385992,cycle)
    `expect("io_rd",io_rd,926385992,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5638024;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,1229940353,cycle)
    `expect("io_rd",io_rd,1229940353,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd4921606;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,1047364631,cycle)
    `expect("io_rd",io_rd,1047364631,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3968110;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,1087702566,cycle)
    `expect("io_rd",io_rd,1087702566,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd6043337;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,1066495931,cycle)
    `expect("io_rd",io_rd,1066495931,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd4532835;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,1030708799,cycle)
    `expect("io_rd",io_rd,1030708799,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd4707598;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,1108948742,cycle)
    `expect("io_rd",io_rd,1108948742,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1978477;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,919231710,cycle)
    `expect("io_rd",io_rd,919231710,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3377973;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,974269428,cycle)
    `expect("io_rd",io_rd,974269428,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2099837;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,672874995,cycle)
    `expect("io_rd",io_rd,672874995,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd6432280;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,843899143,cycle)
    `expect("io_rd",io_rd,843899143,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd4782390;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,686800673,cycle)
    `expect("io_rd",io_rd,686800673,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 19'd291799;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,822921814,cycle)
    `expect("io_rd",io_rd,822921814,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 17'd84247;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,721724006,cycle)
    `expect("io_rd",io_rd,721724006,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2346101;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,577506467,cycle)
    `expect("io_rd",io_rd,577506467,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3369252;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,399230887,cycle)
    `expect("io_rd",io_rd,399230887,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2133625;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,346077284,cycle)
    `expect("io_rd",io_rd,346077284,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3627415;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,546466083,cycle)
    `expect("io_rd",io_rd,546466083,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd2020252;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,542251100,cycle)
    `expect("io_rd",io_rd,542251100,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 19'd368157;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,559425476,cycle)
    `expect("io_rd",io_rd,559425476,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2261868;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,489301862,cycle)
    `expect("io_rd",io_rd,489301862,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 20'd608904;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,323311033,cycle)
    `expect("io_rd",io_rd,323311033,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2976283;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,411626825,cycle)
    `expect("io_rd",io_rd,411626825,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1337586;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,256695823,cycle)
    `expect("io_rd",io_rd,256695823,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5592101;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,608546810,cycle)
    `expect("io_rd",io_rd,608546810,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3350711;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,479785939,cycle)
    `expect("io_rd",io_rd,479785939,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd4087275;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,844184471,cycle)
    `expect("io_rd",io_rd,844184471,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 20'd842209;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,640125318,cycle)
    `expect("io_rd",io_rd,640125318,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5544299;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,931753912,cycle)
    `expect("io_rd",io_rd,931753912,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3736874;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,614390990,cycle)
    `expect("io_rd",io_rd,614390990,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd4981660;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,911860593,cycle)
    `expect("io_rd",io_rd,911860593,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1242097;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,679588111,cycle)
    `expect("io_rd",io_rd,679588111,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3488486;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,936282165,cycle)
    `expect("io_rd",io_rd,936282165,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3621113;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,657096477,cycle)
    `expect("io_rd",io_rd,657096477,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5754850;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,833258297,cycle)
    `expect("io_rd",io_rd,833258297,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1864866;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,646995140,cycle)
    `expect("io_rd",io_rd,646995140,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2896942;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,892020136,cycle)
    `expect("io_rd",io_rd,892020136,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5333414;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,792366990,cycle)
    `expect("io_rd",io_rd,792366990,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1643584;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,701093171,cycle)
    `expect("io_rd",io_rd,701093171,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5909719;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,884140859,cycle)
    `expect("io_rd",io_rd,884140859,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3996320;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,723442639,cycle)
    `expect("io_rd",io_rd,723442639,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 19'd271852;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,832420644,cycle)
    `expect("io_rd",io_rd,832420644,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 20'd642436;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,643323415,cycle)
    `expect("io_rd",io_rd,643323415,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2552739;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,541631484,cycle)
    `expect("io_rd",io_rd,541631484,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 19'd524105;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,294394204,cycle)
    `expect("io_rd",io_rd,294394204,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5132214;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,459759565,cycle)
    `expect("io_rd",io_rd,459759565,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd4702834;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,449286181,cycle)
    `expect("io_rd",io_rd,449286181,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd2096459;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,698733208,cycle)
    `expect("io_rd",io_rd,698733208,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5430981;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,851950742,cycle)
    `expect("io_rd",io_rd,851950742,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2264160;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,748769705,cycle)
    `expect("io_rd",io_rd,748769705,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3907476;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,907655057,cycle)
    `expect("io_rd",io_rd,907655057,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 19'd467117;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,561645029,cycle)
    `expect("io_rd",io_rd,561645029,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 19'd371410;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,647259457,cycle)
    `expect("io_rd",io_rd,647259457,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd4964927;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,495823467,cycle)
    `expect("io_rd",io_rd,495823467,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd6317945;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,558737257,cycle)
    `expect("io_rd",io_rd,558737257,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1289457;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,585516908,cycle)
    `expect("io_rd",io_rd,585516908,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2243445;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,819980469,cycle)
    `expect("io_rd",io_rd,819980469,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3586594;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,741631080,cycle)
    `expect("io_rd",io_rd,741631080,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1663467;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,622448360,cycle)
    `expect("io_rd",io_rd,622448360,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5622155;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,685468812,cycle)
    `expect("io_rd",io_rd,685468812,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3134711;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,589373306,cycle)
    `expect("io_rd",io_rd,589373306,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2678331;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,822543978,cycle)
    `expect("io_rd",io_rd,822543978,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd2059659;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,664856218,cycle)
    `expect("io_rd",io_rd,664856218,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd4484156;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,790163859,cycle)
    `expect("io_rd",io_rd,790163859,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5059035;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,683942740,cycle)
    `expect("io_rd",io_rd,683942740,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5785310;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,871761733,cycle)
    `expect("io_rd",io_rd,871761733,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 20'd967456;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,796270924,cycle)
    `expect("io_rd",io_rd,796270924,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1492271;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,918206011,cycle)
    `expect("io_rd",io_rd,918206011,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd6224114;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,796760640,cycle)
    `expect("io_rd",io_rd,796760640,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1784162;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,578020491,cycle)
    `expect("io_rd",io_rd,578020491,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd4076917;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,788402304,cycle)
    `expect("io_rd",io_rd,788402304,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3879170;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,673851527,cycle)
    `expect("io_rd",io_rd,673851527,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3603745;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,867692375,cycle)
    `expect("io_rd",io_rd,867692375,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd4216693;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,774381708,cycle)
    `expect("io_rd",io_rd,774381708,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3928363;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,840003025,cycle)
    `expect("io_rd",io_rd,840003025,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3110146;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,830401008,cycle)
    `expect("io_rd",io_rd,830401008,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1624862;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,744089193,cycle)
    `expect("io_rd",io_rd,744089193,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5232199;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,819370747,cycle)
    `expect("io_rd",io_rd,819370747,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2273772;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,596509781,cycle)
    `expect("io_rd",io_rd,596509781,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2751468;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,758761978,cycle)
    `expect("io_rd",io_rd,758761978,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 19'd509547;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,517095859,cycle)
    `expect("io_rd",io_rd,517095859,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 19'd265745;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,544521441,cycle)
    `expect("io_rd",io_rd,544521441,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd6101946;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,500510861,cycle)
    `expect("io_rd",io_rd,500510861,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3031531;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,385792560,cycle)
    `expect("io_rd",io_rd,385792560,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 19'd491313;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,584026485,cycle)
    `expect("io_rd",io_rd,584026485,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5274800;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,713206152,cycle)
    `expect("io_rd",io_rd,713206152,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3605440;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,651898760,cycle)
    `expect("io_rd",io_rd,651898760,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd6518463;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,894361079,cycle)
    `expect("io_rd",io_rd,894361079,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5071680;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,829413159,cycle)
    `expect("io_rd",io_rd,829413159,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd2093630;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,1047576927,cycle)
    `expect("io_rd",io_rd,1047576927,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5398988;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,1062905776,cycle)
    `expect("io_rd",io_rd,1062905776,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5242265;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,944577786,cycle)
    `expect("io_rd",io_rd,944577786,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd6433389;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,1076021474,cycle)
    `expect("io_rd",io_rd,1076021474,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2235905;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,911170107,cycle)
    `expect("io_rd",io_rd,911170107,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5611285;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,1207725824,cycle)
    `expect("io_rd",io_rd,1207725824,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 16'd54395;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,742228124,cycle)
    `expect("io_rd",io_rd,742228124,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5138119;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,1014009433,cycle)
    `expect("io_rd",io_rd,1014009433,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1520973;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,465079082,cycle)
    `expect("io_rd",io_rd,465079082,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1314115;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,723587200,cycle)
    `expect("io_rd",io_rd,723587200,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd4561293;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,532350895,cycle)
    `expect("io_rd",io_rd,532350895,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1362115;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,512409389,cycle)
    `expect("io_rd",io_rd,512409389,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd4466288;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,682945354,cycle)
    `expect("io_rd",io_rd,682945354,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3432122;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,556931905,cycle)
    `expect("io_rd",io_rd,556931905,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 16'd62840;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,657108315,cycle)
    `expect("io_rd",io_rd,657108315,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd6460228;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,769941016,cycle)
    `expect("io_rd",io_rd,769941016,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5437517;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,660982780,cycle)
    `expect("io_rd",io_rd,660982780,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd6401057;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,1014155774,cycle)
    `expect("io_rd",io_rd,1014155774,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5131892;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,1001920904,cycle)
    `expect("io_rd",io_rd,1001920904,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3236035;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,1207505894,cycle)
    `expect("io_rd",io_rd,1207505894,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2682061;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,1046529314,cycle)
    `expect("io_rd",io_rd,1046529314,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5072870;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,978969875,cycle)
    `expect("io_rd",io_rd,978969875,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2820710;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,755407874,cycle)
    `expect("io_rd",io_rd,755407874,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd6094390;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,940671253,cycle)
    `expect("io_rd",io_rd,940671253,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2759138;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,748688190,cycle)
    `expect("io_rd",io_rd,748688190,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5628923;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,1083446954,cycle)
    `expect("io_rd",io_rd,1083446954,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3151706;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,797557819,cycle)
    `expect("io_rd",io_rd,797557819,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5789510;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,1100759344,cycle)
    `expect("io_rd",io_rd,1100759344,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2155448;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,769179687,cycle)
    `expect("io_rd",io_rd,769179687,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2874721;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,970796282,cycle)
    `expect("io_rd",io_rd,970796282,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 19'd281161;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,586173089,cycle)
    `expect("io_rd",io_rd,586173089,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3481221;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,703107056,cycle)
    `expect("io_rd",io_rd,703107056,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2986808;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,406986845,cycle)
    `expect("io_rd",io_rd,406986845,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3983720;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,622426425,cycle)
    `expect("io_rd",io_rd,622426425,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 19'd412983;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,465913700,cycle)
    `expect("io_rd",io_rd,465913700,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1063095;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,626878998,cycle)
    `expect("io_rd",io_rd,626878998,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1622002;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,397504162,cycle)
    `expect("io_rd",io_rd,397504162,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5250644;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,513424843,cycle)
    `expect("io_rd",io_rd,513424843,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5490817;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,503428014,cycle)
    `expect("io_rd",io_rd,503428014,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd4227365;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,789665489,cycle)
    `expect("io_rd",io_rd,789665489,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 19'd265325;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,785860607,cycle)
    `expect("io_rd",io_rd,785860607,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5444103;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,997043021,cycle)
    `expect("io_rd",io_rd,997043021,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2898025;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,627905187,cycle)
    `expect("io_rd",io_rd,627905187,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5575401;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,898149350,cycle)
    `expect("io_rd",io_rd,898149350,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3307685;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,681350137,cycle)
    `expect("io_rd",io_rd,681350137,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1550827;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,900734250,cycle)
    `expect("io_rd",io_rd,900734250,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd4526291;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,812287173,cycle)
    `expect("io_rd",io_rd,812287173,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 20'd984471;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,602092453,cycle)
    `expect("io_rd",io_rd,602092453,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5050796;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,782531321,cycle)
    `expect("io_rd",io_rd,782531321,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2729143;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,516429130,cycle)
    `expect("io_rd",io_rd,516429130,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5478033;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,900598525,cycle)
    `expect("io_rd",io_rd,900598525,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3993437;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,710064824,cycle)
    `expect("io_rd",io_rd,710064824,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3266401;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,952971437,cycle)
    `expect("io_rd",io_rd,952971437,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5750242;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,935364478,cycle)
    `expect("io_rd",io_rd,935364478,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2222211;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,831773044,cycle)
    `expect("io_rd",io_rd,831773044,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5195948;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,1000966519,cycle)
    `expect("io_rd",io_rd,1000966519,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3748669;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,778292562,cycle)
    `expect("io_rd",io_rd,778292562,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1235145;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,851986343,cycle)
    `expect("io_rd",io_rd,851986343,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5856371;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,853935527,cycle)
    `expect("io_rd",io_rd,853935527,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3281633;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,696338836,cycle)
    `expect("io_rd",io_rd,696338836,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2309787;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,818441188,cycle)
    `expect("io_rd",io_rd,818441188,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 19'd484145;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,595620748,cycle)
    `expect("io_rd",io_rd,595620748,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 20'd879764;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,600031496,cycle)
    `expect("io_rd",io_rd,600031496,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5523706;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,510240146,cycle)
    `expect("io_rd",io_rd,510240146,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1858530;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,355978669,cycle)
    `expect("io_rd",io_rd,355978669,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1384884;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,578462621,cycle)
    `expect("io_rd",io_rd,578462621,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3761228;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,576481505,cycle)
    `expect("io_rd",io_rd,576481505,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5266540;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,696225050,cycle)
    `expect("io_rd",io_rd,696225050,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1990266;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,599815121,cycle)
    `expect("io_rd",io_rd,599815121,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5626106;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,886050674,cycle)
    `expect("io_rd",io_rd,886050674,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd4898329;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,817326024,cycle)
    `expect("io_rd",io_rd,817326024,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3691872;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,978220274,cycle)
    `expect("io_rd",io_rd,978220274,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5163455;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,963994882,cycle)
    `expect("io_rd",io_rd,963994882,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3011076;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,929346102,cycle)
    `expect("io_rd",io_rd,929346102,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 19'd279086;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,817978377,cycle)
    `expect("io_rd",io_rd,817978377,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd6386225;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,862389660,cycle)
    `expect("io_rd",io_rd,862389660,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2277539;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,558376401,cycle)
    `expect("io_rd",io_rd,558376401,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd6367972;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,944149436,cycle)
    `expect("io_rd",io_rd,944149436,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3376834;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,685673529,cycle)
    `expect("io_rd",io_rd,685673529,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3930896;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,1079138001,cycle)
    `expect("io_rd",io_rd,1079138001,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd3888914;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,835867777,cycle)
    `expect("io_rd",io_rd,835867777,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1527081;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,837427649,cycle)
    `expect("io_rd",io_rd,837427649,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 20'd860402;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,661827168,cycle)
    `expect("io_rd",io_rd,661827168,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5988525;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,699675041,cycle)
    `expect("io_rd",io_rd,699675041,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1139955;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,439158707,cycle)
    `expect("io_rd",io_rd,439158707,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 21'd1719560;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,660047003,cycle)
    `expect("io_rd",io_rd,660047003,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2545807;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,492069484,cycle)
    `expect("io_rd",io_rd,492069484,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd4320630;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,654537700,cycle)
    `expect("io_rd",io_rd,654537700,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5972233;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,636459697,cycle)
    `expect("io_rd",io_rd,636459697,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5164239;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,826831568,cycle)
    `expect("io_rd",io_rd,826831568,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2904887;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,952508488,cycle)
    `expect("io_rd",io_rd,952508488,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 23'd5956804;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,1116178979,cycle)
    `expect("io_rd",io_rd,1116178979,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2955722;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,903301560,cycle)
    `expect("io_rd",io_rd,903301560,cycle)
    io_valid = 1'd0;
    io_valid = 1'd1;
    io_insn = 6'd43;
    io_rs1 = 22'd2864281;
    #(1*`CLK_PERIOD)     io_valid = 1'd0;
    #(1*`CLK_PERIOD)     io_valid = 1'd1;
    io_insn = 6'd59;
    #(1*`CLK_PERIOD)     `expect("io_rd",io_rd,967967175,cycle)
    `expect("io_rd",io_rd,967967175,cycle)
    io_valid = 1'd0;

    #`CLK_PERIOD $display("\t **Ran through all test vectors**"); $finish;

  end
endmodule