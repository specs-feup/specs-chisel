module SCIEPipelined #(parameter XLEN = 32)(
  input         clock,
  input         reset,
  input         valid,
  input  [31:0] insn,
  input  [31:0] rs1,
  input  [31:0] rs2,
  output [31:0] rd
);
  reg [31:0] coeffs_0;
  reg [31:0] coeffs_1;
  reg [31:0] coeffs_2;
  reg [31:0] coeffs_3;
  reg [31:0] coeffs_4;
  reg [31:0] coeffs_5;
  reg [31:0] coeffs_6;
  reg [31:0] coeffs_7;
  reg [31:0] coeffs_8;
  reg [31:0] coeffs_9;
  reg [31:0] coeffs_10;
  reg [31:0] coeffs_11;
  reg [31:0] coeffs_12;
  reg [31:0] coeffs_13;
  reg [31:0] coeffs_14;
  reg [31:0] coeffs_15;
  reg [31:0] coeffs_16;
  reg [31:0] coeffs_17;
  reg [31:0] coeffs_18;
  reg [31:0] coeffs_19;
  reg [31:0] coeffs_20;
  reg [31:0] coeffs_21;
  reg [31:0] coeffs_22;
  reg [31:0] coeffs_23;
  reg [31:0] coeffs_24;
  reg [31:0] coeffs_25;
  reg [31:0] coeffs_26;
  reg [31:0] coeffs_27;
  reg [31:0] coeffs_28;
  reg [31:0] coeffs_29;
  reg [31:0] coeffs_30;
  reg [31:0] coeffs_31;
  reg [31:0] coeffs_32;
  reg [31:0] coeffs_33;
  reg [31:0] coeffs_34;
  reg [31:0] coeffs_35;
  reg [31:0] coeffs_36;
  reg [31:0] coeffs_37;
  reg [31:0] coeffs_38;
  reg [31:0] coeffs_39;
  reg [31:0] coeffs_40;
  reg [31:0] coeffs_41;
  reg [31:0] coeffs_42;
  reg [31:0] coeffs_43;
  reg [31:0] coeffs_44;
  reg [31:0] coeffs_45;
  reg [31:0] coeffs_46;
  reg [31:0] coeffs_47;
  reg [31:0] coeffs_48;
  reg [31:0] coeffs_49;
  reg [31:0] coeffs_50;
  reg [31:0] coeffs_51;
  reg [31:0] coeffs_52;
  reg [31:0] coeffs_53;
  reg [31:0] coeffs_54;
  reg [31:0] coeffs_55;
  reg [31:0] coeffs_56;
  reg [31:0] coeffs_57;
  reg [31:0] coeffs_58;
  reg [31:0] coeffs_59;
  reg [31:0] coeffs_60;
  reg [31:0] coeffs_61;
  reg [31:0] coeffs_62;
  reg [31:0] coeffs_63;
  reg [31:0] coeffs_64;
  reg [31:0] coeffs_65;
  reg [31:0] coeffs_66;
  reg [31:0] coeffs_67;
  reg [31:0] coeffs_68;
  reg [31:0] coeffs_69;
  reg [31:0] coeffs_70;
  reg [31:0] coeffs_71;
  reg [31:0] coeffs_72;
  reg [31:0] coeffs_73;
  reg [31:0] coeffs_74;
  reg [31:0] coeffs_75;
  reg [31:0] coeffs_76;
  reg [31:0] coeffs_77;
  reg [31:0] coeffs_78;
  reg [31:0] coeffs_79;
  reg [31:0] coeffs_80;
  reg [31:0] coeffs_81;
  reg [31:0] coeffs_82;
  reg [31:0] coeffs_83;
  reg [31:0] coeffs_84;
  reg [31:0] coeffs_85;
  reg [31:0] coeffs_86;
  reg [31:0] coeffs_87;
  reg [31:0] coeffs_88;
  reg [31:0] coeffs_89;
  reg [31:0] coeffs_90;
  reg [31:0] coeffs_91;
  reg [31:0] coeffs_92;
  reg [31:0] coeffs_93;
  reg [31:0] coeffs_94;
  reg [31:0] coeffs_95;
  reg [31:0] coeffs_96;
  reg [31:0] coeffs_97;
  reg [31:0] coeffs_98;
  reg [31:0] coeffs_99;
  reg [31:0] data_0;
  reg [31:0] data_1;
  reg [31:0] data_2;
  reg [31:0] data_3;
  reg [31:0] data_4;
  reg [31:0] data_5;
  reg [31:0] data_6;
  reg [31:0] data_7;
  reg [31:0] data_8;
  reg [31:0] data_9;
  reg [31:0] data_10;
  reg [31:0] data_11;
  reg [31:0] data_12;
  reg [31:0] data_13;
  reg [31:0] data_14;
  reg [31:0] data_15;
  reg [31:0] data_16;
  reg [31:0] data_17;
  reg [31:0] data_18;
  reg [31:0] data_19;
  reg [31:0] data_20;
  reg [31:0] data_21;
  reg [31:0] data_22;
  reg [31:0] data_23;
  reg [31:0] data_24;
  reg [31:0] data_25;
  reg [31:0] data_26;
  reg [31:0] data_27;
  reg [31:0] data_28;
  reg [31:0] data_29;
  reg [31:0] data_30;
  reg [31:0] data_31;
  reg [31:0] data_32;
  reg [31:0] data_33;
  reg [31:0] data_34;
  reg [31:0] data_35;
  reg [31:0] data_36;
  reg [31:0] data_37;
  reg [31:0] data_38;
  reg [31:0] data_39;
  reg [31:0] data_40;
  reg [31:0] data_41;
  reg [31:0] data_42;
  reg [31:0] data_43;
  reg [31:0] data_44;
  reg [31:0] data_45;
  reg [31:0] data_46;
  reg [31:0] data_47;
  reg [31:0] data_48;
  reg [31:0] data_49;
  reg [31:0] data_50;
  reg [31:0] data_51;
  reg [31:0] data_52;
  reg [31:0] data_53;
  reg [31:0] data_54;
  reg [31:0] data_55;
  reg [31:0] data_56;
  reg [31:0] data_57;
  reg [31:0] data_58;
  reg [31:0] data_59;
  reg [31:0] data_60;
  reg [31:0] data_61;
  reg [31:0] data_62;
  reg [31:0] data_63;
  reg [31:0] data_64;
  reg [31:0] data_65;
  reg [31:0] data_66;
  reg [31:0] data_67;
  reg [31:0] data_68;
  reg [31:0] data_69;
  reg [31:0] data_70;
  reg [31:0] data_71;
  reg [31:0] data_72;
  reg [31:0] data_73;
  reg [31:0] data_74;
  reg [31:0] data_75;
  reg [31:0] data_76;
  reg [31:0] data_77;
  reg [31:0] data_78;
  reg [31:0] data_79;
  reg [31:0] data_80;
  reg [31:0] data_81;
  reg [31:0] data_82;
  reg [31:0] data_83;
  reg [31:0] data_84;
  reg [31:0] data_85;
  reg [31:0] data_86;
  reg [31:0] data_87;
  reg [31:0] data_88;
  reg [31:0] data_89;
  reg [31:0] data_90;
  reg [31:0] data_91;
  reg [31:0] data_92;
  reg [31:0] data_93;
  reg [31:0] data_94;
  reg [31:0] data_95;
  reg [31:0] data_96;
  reg [31:0] data_97;
  reg [31:0] data_98;
  reg [31:0] data_99;
  reg [63:0] result;
  wire [31:0] _GEN_101 = 7'h1 == rs2[6:0] ? coeffs_1 : coeffs_0;
  wire [31:0] _GEN_102 = 7'h2 == rs2[6:0] ? coeffs_2 : _GEN_101;
  wire [31:0] _GEN_103 = 7'h3 == rs2[6:0] ? coeffs_3 : _GEN_102;
  wire [31:0] _GEN_104 = 7'h4 == rs2[6:0] ? coeffs_4 : _GEN_103;
  wire [31:0] _GEN_105 = 7'h5 == rs2[6:0] ? coeffs_5 : _GEN_104;
  wire [31:0] _GEN_106 = 7'h6 == rs2[6:0] ? coeffs_6 : _GEN_105;
  wire [31:0] _GEN_107 = 7'h7 == rs2[6:0] ? coeffs_7 : _GEN_106;
  wire [31:0] _GEN_108 = 7'h8 == rs2[6:0] ? coeffs_8 : _GEN_107;
  wire [31:0] _GEN_109 = 7'h9 == rs2[6:0] ? coeffs_9 : _GEN_108;
  wire [31:0] _GEN_110 = 7'ha == rs2[6:0] ? coeffs_10 : _GEN_109;
  wire [31:0] _GEN_111 = 7'hb == rs2[6:0] ? coeffs_11 : _GEN_110;
  wire [31:0] _GEN_112 = 7'hc == rs2[6:0] ? coeffs_12 : _GEN_111;
  wire [31:0] _GEN_113 = 7'hd == rs2[6:0] ? coeffs_13 : _GEN_112;
  wire [31:0] _GEN_114 = 7'he == rs2[6:0] ? coeffs_14 : _GEN_113;
  wire [31:0] _GEN_115 = 7'hf == rs2[6:0] ? coeffs_15 : _GEN_114;
  wire [31:0] _GEN_116 = 7'h10 == rs2[6:0] ? coeffs_16 : _GEN_115;
  wire [31:0] _GEN_117 = 7'h11 == rs2[6:0] ? coeffs_17 : _GEN_116;
  wire [31:0] _GEN_118 = 7'h12 == rs2[6:0] ? coeffs_18 : _GEN_117;
  wire [31:0] _GEN_119 = 7'h13 == rs2[6:0] ? coeffs_19 : _GEN_118;
  wire [31:0] _GEN_120 = 7'h14 == rs2[6:0] ? coeffs_20 : _GEN_119;
  wire [31:0] _GEN_121 = 7'h15 == rs2[6:0] ? coeffs_21 : _GEN_120;
  wire [31:0] _GEN_122 = 7'h16 == rs2[6:0] ? coeffs_22 : _GEN_121;
  wire [31:0] _GEN_123 = 7'h17 == rs2[6:0] ? coeffs_23 : _GEN_122;
  wire [31:0] _GEN_124 = 7'h18 == rs2[6:0] ? coeffs_24 : _GEN_123;
  wire [31:0] _GEN_125 = 7'h19 == rs2[6:0] ? coeffs_25 : _GEN_124;
  wire [31:0] _GEN_126 = 7'h1a == rs2[6:0] ? coeffs_26 : _GEN_125;
  wire [31:0] _GEN_127 = 7'h1b == rs2[6:0] ? coeffs_27 : _GEN_126;
  wire [31:0] _GEN_128 = 7'h1c == rs2[6:0] ? coeffs_28 : _GEN_127;
  wire [31:0] _GEN_129 = 7'h1d == rs2[6:0] ? coeffs_29 : _GEN_128;
  wire [31:0] _GEN_130 = 7'h1e == rs2[6:0] ? coeffs_30 : _GEN_129;
  wire [31:0] _GEN_131 = 7'h1f == rs2[6:0] ? coeffs_31 : _GEN_130;
  wire [31:0] _GEN_132 = 7'h20 == rs2[6:0] ? coeffs_32 : _GEN_131;
  wire [31:0] _GEN_133 = 7'h21 == rs2[6:0] ? coeffs_33 : _GEN_132;
  wire [31:0] _GEN_134 = 7'h22 == rs2[6:0] ? coeffs_34 : _GEN_133;
  wire [31:0] _GEN_135 = 7'h23 == rs2[6:0] ? coeffs_35 : _GEN_134;
  wire [31:0] _GEN_136 = 7'h24 == rs2[6:0] ? coeffs_36 : _GEN_135;
  wire [31:0] _GEN_137 = 7'h25 == rs2[6:0] ? coeffs_37 : _GEN_136;
  wire [31:0] _GEN_138 = 7'h26 == rs2[6:0] ? coeffs_38 : _GEN_137;
  wire [31:0] _GEN_139 = 7'h27 == rs2[6:0] ? coeffs_39 : _GEN_138;
  wire [31:0] _GEN_140 = 7'h28 == rs2[6:0] ? coeffs_40 : _GEN_139;
  wire [31:0] _GEN_141 = 7'h29 == rs2[6:0] ? coeffs_41 : _GEN_140;
  wire [31:0] _GEN_142 = 7'h2a == rs2[6:0] ? coeffs_42 : _GEN_141;
  wire [31:0] _GEN_143 = 7'h2b == rs2[6:0] ? coeffs_43 : _GEN_142;
  wire [31:0] _GEN_144 = 7'h2c == rs2[6:0] ? coeffs_44 : _GEN_143;
  wire [31:0] _GEN_145 = 7'h2d == rs2[6:0] ? coeffs_45 : _GEN_144;
  wire [31:0] _GEN_146 = 7'h2e == rs2[6:0] ? coeffs_46 : _GEN_145;
  wire [31:0] _GEN_147 = 7'h2f == rs2[6:0] ? coeffs_47 : _GEN_146;
  wire [31:0] _GEN_148 = 7'h30 == rs2[6:0] ? coeffs_48 : _GEN_147;
  wire [31:0] _GEN_149 = 7'h31 == rs2[6:0] ? coeffs_49 : _GEN_148;
  wire [31:0] _GEN_150 = 7'h32 == rs2[6:0] ? coeffs_50 : _GEN_149;
  wire [31:0] _GEN_151 = 7'h33 == rs2[6:0] ? coeffs_51 : _GEN_150;
  wire [31:0] _GEN_152 = 7'h34 == rs2[6:0] ? coeffs_52 : _GEN_151;
  wire [31:0] _GEN_153 = 7'h35 == rs2[6:0] ? coeffs_53 : _GEN_152;
  wire [31:0] _GEN_154 = 7'h36 == rs2[6:0] ? coeffs_54 : _GEN_153;
  wire [31:0] _GEN_155 = 7'h37 == rs2[6:0] ? coeffs_55 : _GEN_154;
  wire [31:0] _GEN_156 = 7'h38 == rs2[6:0] ? coeffs_56 : _GEN_155;
  wire [31:0] _GEN_157 = 7'h39 == rs2[6:0] ? coeffs_57 : _GEN_156;
  wire [31:0] _GEN_158 = 7'h3a == rs2[6:0] ? coeffs_58 : _GEN_157;
  wire [31:0] _GEN_159 = 7'h3b == rs2[6:0] ? coeffs_59 : _GEN_158;
  wire [31:0] _GEN_160 = 7'h3c == rs2[6:0] ? coeffs_60 : _GEN_159;
  wire [31:0] _GEN_161 = 7'h3d == rs2[6:0] ? coeffs_61 : _GEN_160;
  wire [31:0] _GEN_162 = 7'h3e == rs2[6:0] ? coeffs_62 : _GEN_161;
  wire [31:0] _GEN_163 = 7'h3f == rs2[6:0] ? coeffs_63 : _GEN_162;
  wire [31:0] _GEN_164 = 7'h40 == rs2[6:0] ? coeffs_64 : _GEN_163;
  wire [31:0] _GEN_165 = 7'h41 == rs2[6:0] ? coeffs_65 : _GEN_164;
  wire [31:0] _GEN_166 = 7'h42 == rs2[6:0] ? coeffs_66 : _GEN_165;
  wire [31:0] _GEN_167 = 7'h43 == rs2[6:0] ? coeffs_67 : _GEN_166;
  wire [31:0] _GEN_168 = 7'h44 == rs2[6:0] ? coeffs_68 : _GEN_167;
  wire [31:0] _GEN_169 = 7'h45 == rs2[6:0] ? coeffs_69 : _GEN_168;
  wire [31:0] _GEN_170 = 7'h46 == rs2[6:0] ? coeffs_70 : _GEN_169;
  wire [31:0] _GEN_171 = 7'h47 == rs2[6:0] ? coeffs_71 : _GEN_170;
  wire [31:0] _GEN_172 = 7'h48 == rs2[6:0] ? coeffs_72 : _GEN_171;
  wire [31:0] _GEN_173 = 7'h49 == rs2[6:0] ? coeffs_73 : _GEN_172;
  wire [31:0] _GEN_174 = 7'h4a == rs2[6:0] ? coeffs_74 : _GEN_173;
  wire [31:0] _GEN_175 = 7'h4b == rs2[6:0] ? coeffs_75 : _GEN_174;
  wire [31:0] _GEN_176 = 7'h4c == rs2[6:0] ? coeffs_76 : _GEN_175;
  wire [31:0] _GEN_177 = 7'h4d == rs2[6:0] ? coeffs_77 : _GEN_176;
  wire [31:0] _GEN_178 = 7'h4e == rs2[6:0] ? coeffs_78 : _GEN_177;
  wire [31:0] _GEN_179 = 7'h4f == rs2[6:0] ? coeffs_79 : _GEN_178;
  wire [31:0] _GEN_180 = 7'h50 == rs2[6:0] ? coeffs_80 : _GEN_179;
  wire [31:0] _GEN_181 = 7'h51 == rs2[6:0] ? coeffs_81 : _GEN_180;
  wire [31:0] _GEN_182 = 7'h52 == rs2[6:0] ? coeffs_82 : _GEN_181;
  wire [31:0] _GEN_183 = 7'h53 == rs2[6:0] ? coeffs_83 : _GEN_182;
  wire [31:0] _GEN_184 = 7'h54 == rs2[6:0] ? coeffs_84 : _GEN_183;
  wire [31:0] _GEN_185 = 7'h55 == rs2[6:0] ? coeffs_85 : _GEN_184;
  wire [31:0] _GEN_186 = 7'h56 == rs2[6:0] ? coeffs_86 : _GEN_185;
  wire [31:0] _GEN_187 = 7'h57 == rs2[6:0] ? coeffs_87 : _GEN_186;
  wire [31:0] _GEN_188 = 7'h58 == rs2[6:0] ? coeffs_88 : _GEN_187;
  wire [31:0] _GEN_189 = 7'h59 == rs2[6:0] ? coeffs_89 : _GEN_188;
  wire [31:0] _GEN_190 = 7'h5a == rs2[6:0] ? coeffs_90 : _GEN_189;
  wire [31:0] _GEN_191 = 7'h5b == rs2[6:0] ? coeffs_91 : _GEN_190;
  wire [31:0] _GEN_192 = 7'h5c == rs2[6:0] ? coeffs_92 : _GEN_191;
  wire [31:0] _GEN_193 = 7'h5d == rs2[6:0] ? coeffs_93 : _GEN_192;
  wire [31:0] _GEN_194 = 7'h5e == rs2[6:0] ? coeffs_94 : _GEN_193;
  wire [31:0] _GEN_195 = 7'h5f == rs2[6:0] ? coeffs_95 : _GEN_194;
  wire [31:0] _GEN_196 = 7'h60 == rs2[6:0] ? coeffs_96 : _GEN_195;
  wire [31:0] _GEN_197 = 7'h61 == rs2[6:0] ? coeffs_97 : _GEN_196;
  wire [31:0] _GEN_198 = 7'h62 == rs2[6:0] ? coeffs_98 : _GEN_197;
  wire [31:0] _GEN_199 = 7'h63 == rs2[6:0] ? coeffs_99 : _GEN_198;
  wire [63:0] _result_T_1 = data_0 * coeffs_0;
  wire [63:0] _result_T_2 = data_1 * coeffs_1;
  wire [63:0] _result_T_3 = data_2 * coeffs_2;
  wire [63:0] _result_T_4 = data_3 * coeffs_3;
  wire [63:0] _result_T_5 = data_4 * coeffs_4;
  wire [63:0] _result_T_6 = data_5 * coeffs_5;
  wire [63:0] _result_T_7 = data_6 * coeffs_6;
  wire [63:0] _result_T_8 = data_7 * coeffs_7;
  wire [63:0] _result_T_9 = data_8 * coeffs_8;
  wire [63:0] _result_T_10 = data_9 * coeffs_9;
  wire [63:0] _result_T_11 = data_10 * coeffs_10;
  wire [63:0] _result_T_12 = data_11 * coeffs_11;
  wire [63:0] _result_T_13 = data_12 * coeffs_12;
  wire [63:0] _result_T_14 = data_13 * coeffs_13;
  wire [63:0] _result_T_15 = data_14 * coeffs_14;
  wire [63:0] _result_T_16 = data_15 * coeffs_15;
  wire [63:0] _result_T_17 = data_16 * coeffs_16;
  wire [63:0] _result_T_18 = data_17 * coeffs_17;
  wire [63:0] _result_T_19 = data_18 * coeffs_18;
  wire [63:0] _result_T_20 = data_19 * coeffs_19;
  wire [63:0] _result_T_21 = data_20 * coeffs_20;
  wire [63:0] _result_T_22 = data_21 * coeffs_21;
  wire [63:0] _result_T_23 = data_22 * coeffs_22;
  wire [63:0] _result_T_24 = data_23 * coeffs_23;
  wire [63:0] _result_T_25 = data_24 * coeffs_24;
  wire [63:0] _result_T_26 = data_25 * coeffs_25;
  wire [63:0] _result_T_27 = data_26 * coeffs_26;
  wire [63:0] _result_T_28 = data_27 * coeffs_27;
  wire [63:0] _result_T_29 = data_28 * coeffs_28;
  wire [63:0] _result_T_30 = data_29 * coeffs_29;
  wire [63:0] _result_T_31 = data_30 * coeffs_30;
  wire [63:0] _result_T_32 = data_31 * coeffs_31;
  wire [63:0] _result_T_33 = data_32 * coeffs_32;
  wire [63:0] _result_T_34 = data_33 * coeffs_33;
  wire [63:0] _result_T_35 = data_34 * coeffs_34;
  wire [63:0] _result_T_36 = data_35 * coeffs_35;
  wire [63:0] _result_T_37 = data_36 * coeffs_36;
  wire [63:0] _result_T_38 = data_37 * coeffs_37;
  wire [63:0] _result_T_39 = data_38 * coeffs_38;
  wire [63:0] _result_T_40 = data_39 * coeffs_39;
  wire [63:0] _result_T_41 = data_40 * coeffs_40;
  wire [63:0] _result_T_42 = data_41 * coeffs_41;
  wire [63:0] _result_T_43 = data_42 * coeffs_42;
  wire [63:0] _result_T_44 = data_43 * coeffs_43;
  wire [63:0] _result_T_45 = data_44 * coeffs_44;
  wire [63:0] _result_T_46 = data_45 * coeffs_45;
  wire [63:0] _result_T_47 = data_46 * coeffs_46;
  wire [63:0] _result_T_48 = data_47 * coeffs_47;
  wire [63:0] _result_T_49 = data_48 * coeffs_48;
  wire [63:0] _result_T_50 = data_49 * coeffs_49;
  wire [63:0] _result_T_51 = data_50 * coeffs_50;
  wire [63:0] _result_T_52 = data_51 * coeffs_51;
  wire [63:0] _result_T_53 = data_52 * coeffs_52;
  wire [63:0] _result_T_54 = data_53 * coeffs_53;
  wire [63:0] _result_T_55 = data_54 * coeffs_54;
  wire [63:0] _result_T_56 = data_55 * coeffs_55;
  wire [63:0] _result_T_57 = data_56 * coeffs_56;
  wire [63:0] _result_T_58 = data_57 * coeffs_57;
  wire [63:0] _result_T_59 = data_58 * coeffs_58;
  wire [63:0] _result_T_60 = data_59 * coeffs_59;
  wire [63:0] _result_T_61 = data_60 * coeffs_60;
  wire [63:0] _result_T_62 = data_61 * coeffs_61;
  wire [63:0] _result_T_63 = data_62 * coeffs_62;
  wire [63:0] _result_T_64 = data_63 * coeffs_63;
  wire [63:0] _result_T_65 = data_64 * coeffs_64;
  wire [63:0] _result_T_66 = data_65 * coeffs_65;
  wire [63:0] _result_T_67 = data_66 * coeffs_66;
  wire [63:0] _result_T_68 = data_67 * coeffs_67;
  wire [63:0] _result_T_69 = data_68 * coeffs_68;
  wire [63:0] _result_T_70 = data_69 * coeffs_69;
  wire [63:0] _result_T_71 = data_70 * coeffs_70;
  wire [63:0] _result_T_72 = data_71 * coeffs_71;
  wire [63:0] _result_T_73 = data_72 * coeffs_72;
  wire [63:0] _result_T_74 = data_73 * coeffs_73;
  wire [63:0] _result_T_75 = data_74 * coeffs_74;
  wire [63:0] _result_T_76 = data_75 * coeffs_75;
  wire [63:0] _result_T_77 = data_76 * coeffs_76;
  wire [63:0] _result_T_78 = data_77 * coeffs_77;
  wire [63:0] _result_T_79 = data_78 * coeffs_78;
  wire [63:0] _result_T_80 = data_79 * coeffs_79;
  wire [63:0] _result_T_81 = data_80 * coeffs_80;
  wire [63:0] _result_T_82 = data_81 * coeffs_81;
  wire [63:0] _result_T_83 = data_82 * coeffs_82;
  wire [63:0] _result_T_84 = data_83 * coeffs_83;
  wire [63:0] _result_T_85 = data_84 * coeffs_84;
  wire [63:0] _result_T_86 = data_85 * coeffs_85;
  wire [63:0] _result_T_87 = data_86 * coeffs_86;
  wire [63:0] _result_T_88 = data_87 * coeffs_87;
  wire [63:0] _result_T_89 = data_88 * coeffs_88;
  wire [63:0] _result_T_90 = data_89 * coeffs_89;
  wire [63:0] _result_T_91 = data_90 * coeffs_90;
  wire [63:0] _result_T_92 = data_91 * coeffs_91;
  wire [63:0] _result_T_93 = data_92 * coeffs_92;
  wire [63:0] _result_T_94 = data_93 * coeffs_93;
  wire [63:0] _result_T_95 = data_94 * coeffs_94;
  wire [63:0] _result_T_96 = data_95 * coeffs_95;
  wire [63:0] _result_T_97 = data_96 * coeffs_96;
  wire [63:0] _result_T_98 = data_97 * coeffs_97;
  wire [63:0] _result_T_99 = data_98 * coeffs_98;
  wire [63:0] _result_T_100 = data_99 * coeffs_99;
  wire [63:0] _result_T_102 = _result_T_1 + _result_T_2;
  wire [63:0] _result_T_104 = _result_T_102 + _result_T_3;
  wire [63:0] _result_T_106 = _result_T_104 + _result_T_4;
  wire [63:0] _result_T_108 = _result_T_106 + _result_T_5;
  wire [63:0] _result_T_110 = _result_T_108 + _result_T_6;
  wire [63:0] _result_T_112 = _result_T_110 + _result_T_7;
  wire [63:0] _result_T_114 = _result_T_112 + _result_T_8;
  wire [63:0] _result_T_116 = _result_T_114 + _result_T_9;
  wire [63:0] _result_T_118 = _result_T_116 + _result_T_10;
  wire [63:0] _result_T_120 = _result_T_118 + _result_T_11;
  wire [63:0] _result_T_122 = _result_T_120 + _result_T_12;
  wire [63:0] _result_T_124 = _result_T_122 + _result_T_13;
  wire [63:0] _result_T_126 = _result_T_124 + _result_T_14;
  wire [63:0] _result_T_128 = _result_T_126 + _result_T_15;
  wire [63:0] _result_T_130 = _result_T_128 + _result_T_16;
  wire [63:0] _result_T_132 = _result_T_130 + _result_T_17;
  wire [63:0] _result_T_134 = _result_T_132 + _result_T_18;
  wire [63:0] _result_T_136 = _result_T_134 + _result_T_19;
  wire [63:0] _result_T_138 = _result_T_136 + _result_T_20;
  wire [63:0] _result_T_140 = _result_T_138 + _result_T_21;
  wire [63:0] _result_T_142 = _result_T_140 + _result_T_22;
  wire [63:0] _result_T_144 = _result_T_142 + _result_T_23;
  wire [63:0] _result_T_146 = _result_T_144 + _result_T_24;
  wire [63:0] _result_T_148 = _result_T_146 + _result_T_25;
  wire [63:0] _result_T_150 = _result_T_148 + _result_T_26;
  wire [63:0] _result_T_152 = _result_T_150 + _result_T_27;
  wire [63:0] _result_T_154 = _result_T_152 + _result_T_28;
  wire [63:0] _result_T_156 = _result_T_154 + _result_T_29;
  wire [63:0] _result_T_158 = _result_T_156 + _result_T_30;
  wire [63:0] _result_T_160 = _result_T_158 + _result_T_31;
  wire [63:0] _result_T_162 = _result_T_160 + _result_T_32;
  wire [63:0] _result_T_164 = _result_T_162 + _result_T_33;
  wire [63:0] _result_T_166 = _result_T_164 + _result_T_34;
  wire [63:0] _result_T_168 = _result_T_166 + _result_T_35;
  wire [63:0] _result_T_170 = _result_T_168 + _result_T_36;
  wire [63:0] _result_T_172 = _result_T_170 + _result_T_37;
  wire [63:0] _result_T_174 = _result_T_172 + _result_T_38;
  wire [63:0] _result_T_176 = _result_T_174 + _result_T_39;
  wire [63:0] _result_T_178 = _result_T_176 + _result_T_40;
  wire [63:0] _result_T_180 = _result_T_178 + _result_T_41;
  wire [63:0] _result_T_182 = _result_T_180 + _result_T_42;
  wire [63:0] _result_T_184 = _result_T_182 + _result_T_43;
  wire [63:0] _result_T_186 = _result_T_184 + _result_T_44;
  wire [63:0] _result_T_188 = _result_T_186 + _result_T_45;
  wire [63:0] _result_T_190 = _result_T_188 + _result_T_46;
  wire [63:0] _result_T_192 = _result_T_190 + _result_T_47;
  wire [63:0] _result_T_194 = _result_T_192 + _result_T_48;
  wire [63:0] _result_T_196 = _result_T_194 + _result_T_49;
  wire [63:0] _result_T_198 = _result_T_196 + _result_T_50;
  wire [63:0] _result_T_200 = _result_T_198 + _result_T_51;
  wire [63:0] _result_T_202 = _result_T_200 + _result_T_52;
  wire [63:0] _result_T_204 = _result_T_202 + _result_T_53;
  wire [63:0] _result_T_206 = _result_T_204 + _result_T_54;
  wire [63:0] _result_T_208 = _result_T_206 + _result_T_55;
  wire [63:0] _result_T_210 = _result_T_208 + _result_T_56;
  wire [63:0] _result_T_212 = _result_T_210 + _result_T_57;
  wire [63:0] _result_T_214 = _result_T_212 + _result_T_58;
  wire [63:0] _result_T_216 = _result_T_214 + _result_T_59;
  wire [63:0] _result_T_218 = _result_T_216 + _result_T_60;
  wire [63:0] _result_T_220 = _result_T_218 + _result_T_61;
  wire [63:0] _result_T_222 = _result_T_220 + _result_T_62;
  wire [63:0] _result_T_224 = _result_T_222 + _result_T_63;
  wire [63:0] _result_T_226 = _result_T_224 + _result_T_64;
  wire [63:0] _result_T_228 = _result_T_226 + _result_T_65;
  wire [63:0] _result_T_230 = _result_T_228 + _result_T_66;
  wire [63:0] _result_T_232 = _result_T_230 + _result_T_67;
  wire [63:0] _result_T_234 = _result_T_232 + _result_T_68;
  wire [63:0] _result_T_236 = _result_T_234 + _result_T_69;
  wire [63:0] _result_T_238 = _result_T_236 + _result_T_70;
  wire [63:0] _result_T_240 = _result_T_238 + _result_T_71;
  wire [63:0] _result_T_242 = _result_T_240 + _result_T_72;
  wire [63:0] _result_T_244 = _result_T_242 + _result_T_73;
  wire [63:0] _result_T_246 = _result_T_244 + _result_T_74;
  wire [63:0] _result_T_248 = _result_T_246 + _result_T_75;
  wire [63:0] _result_T_250 = _result_T_248 + _result_T_76;
  wire [63:0] _result_T_252 = _result_T_250 + _result_T_77;
  wire [63:0] _result_T_254 = _result_T_252 + _result_T_78;
  wire [63:0] _result_T_256 = _result_T_254 + _result_T_79;
  wire [63:0] _result_T_258 = _result_T_256 + _result_T_80;
  wire [63:0] _result_T_260 = _result_T_258 + _result_T_81;
  wire [63:0] _result_T_262 = _result_T_260 + _result_T_82;
  wire [63:0] _result_T_264 = _result_T_262 + _result_T_83;
  wire [63:0] _result_T_266 = _result_T_264 + _result_T_84;
  wire [63:0] _result_T_268 = _result_T_266 + _result_T_85;
  wire [63:0] _result_T_270 = _result_T_268 + _result_T_86;
  wire [63:0] _result_T_272 = _result_T_270 + _result_T_87;
  wire [63:0] _result_T_274 = _result_T_272 + _result_T_88;
  wire [63:0] _result_T_276 = _result_T_274 + _result_T_89;
  wire [63:0] _result_T_278 = _result_T_276 + _result_T_90;
  wire [63:0] _result_T_280 = _result_T_278 + _result_T_91;
  wire [63:0] _result_T_282 = _result_T_280 + _result_T_92;
  wire [63:0] _result_T_284 = _result_T_282 + _result_T_93;
  wire [63:0] _result_T_286 = _result_T_284 + _result_T_94;
  wire [63:0] _result_T_288 = _result_T_286 + _result_T_95;
  wire [63:0] _result_T_290 = _result_T_288 + _result_T_96;
  wire [63:0] _result_T_292 = _result_T_290 + _result_T_97;
  wire [63:0] _result_T_294 = _result_T_292 + _result_T_98;
  wire [63:0] _result_T_296 = _result_T_294 + _result_T_99;
  wire [63:0] _result_T_298 = _result_T_296 + _result_T_100;
  wire [63:0] _GEN_200 = insn[6:0] == 7'h3b ? _result_T_298 : result;
  assign rd = result[31:0];
  always @(posedge clock) begin
    if (reset) begin
      coeffs_0 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h0 == rs2[6:0]) begin
          coeffs_0 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_1 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h1 == rs2[6:0]) begin
          coeffs_1 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_2 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h2 == rs2[6:0]) begin
          coeffs_2 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_3 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h3 == rs2[6:0]) begin
          coeffs_3 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_4 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h4 == rs2[6:0]) begin
          coeffs_4 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_5 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h5 == rs2[6:0]) begin
          coeffs_5 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_6 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h6 == rs2[6:0]) begin
          coeffs_6 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_7 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h7 == rs2[6:0]) begin
          coeffs_7 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_8 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h8 == rs2[6:0]) begin
          coeffs_8 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_9 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h9 == rs2[6:0]) begin
          coeffs_9 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_10 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'ha == rs2[6:0]) begin
          coeffs_10 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_11 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'hb == rs2[6:0]) begin
          coeffs_11 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_12 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'hc == rs2[6:0]) begin
          coeffs_12 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_13 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'hd == rs2[6:0]) begin
          coeffs_13 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_14 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'he == rs2[6:0]) begin
          coeffs_14 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_15 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'hf == rs2[6:0]) begin
          coeffs_15 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_16 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h10 == rs2[6:0]) begin
          coeffs_16 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_17 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h11 == rs2[6:0]) begin
          coeffs_17 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_18 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h12 == rs2[6:0]) begin
          coeffs_18 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_19 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h13 == rs2[6:0]) begin
          coeffs_19 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_20 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h14 == rs2[6:0]) begin
          coeffs_20 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_21 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h15 == rs2[6:0]) begin
          coeffs_21 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_22 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h16 == rs2[6:0]) begin
          coeffs_22 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_23 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h17 == rs2[6:0]) begin
          coeffs_23 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_24 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h18 == rs2[6:0]) begin
          coeffs_24 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_25 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h19 == rs2[6:0]) begin
          coeffs_25 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_26 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h1a == rs2[6:0]) begin
          coeffs_26 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_27 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h1b == rs2[6:0]) begin
          coeffs_27 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_28 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h1c == rs2[6:0]) begin
          coeffs_28 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_29 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h1d == rs2[6:0]) begin
          coeffs_29 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_30 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h1e == rs2[6:0]) begin
          coeffs_30 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_31 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h1f == rs2[6:0]) begin
          coeffs_31 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_32 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h20 == rs2[6:0]) begin
          coeffs_32 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_33 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h21 == rs2[6:0]) begin
          coeffs_33 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_34 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h22 == rs2[6:0]) begin
          coeffs_34 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_35 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h23 == rs2[6:0]) begin
          coeffs_35 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_36 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h24 == rs2[6:0]) begin
          coeffs_36 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_37 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h25 == rs2[6:0]) begin
          coeffs_37 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_38 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h26 == rs2[6:0]) begin
          coeffs_38 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_39 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h27 == rs2[6:0]) begin
          coeffs_39 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_40 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h28 == rs2[6:0]) begin
          coeffs_40 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_41 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h29 == rs2[6:0]) begin
          coeffs_41 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_42 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h2a == rs2[6:0]) begin
          coeffs_42 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_43 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h2b == rs2[6:0]) begin
          coeffs_43 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_44 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h2c == rs2[6:0]) begin
          coeffs_44 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_45 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h2d == rs2[6:0]) begin
          coeffs_45 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_46 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h2e == rs2[6:0]) begin
          coeffs_46 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_47 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h2f == rs2[6:0]) begin
          coeffs_47 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_48 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h30 == rs2[6:0]) begin
          coeffs_48 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_49 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h31 == rs2[6:0]) begin
          coeffs_49 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_50 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h32 == rs2[6:0]) begin
          coeffs_50 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_51 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h33 == rs2[6:0]) begin
          coeffs_51 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_52 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h34 == rs2[6:0]) begin
          coeffs_52 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_53 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h35 == rs2[6:0]) begin
          coeffs_53 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_54 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h36 == rs2[6:0]) begin
          coeffs_54 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_55 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h37 == rs2[6:0]) begin
          coeffs_55 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_56 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h38 == rs2[6:0]) begin
          coeffs_56 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_57 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h39 == rs2[6:0]) begin
          coeffs_57 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_58 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h3a == rs2[6:0]) begin
          coeffs_58 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_59 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h3b == rs2[6:0]) begin
          coeffs_59 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_60 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h3c == rs2[6:0]) begin
          coeffs_60 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_61 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h3d == rs2[6:0]) begin
          coeffs_61 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_62 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h3e == rs2[6:0]) begin
          coeffs_62 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_63 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h3f == rs2[6:0]) begin
          coeffs_63 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_64 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h40 == rs2[6:0]) begin
          coeffs_64 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_65 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h41 == rs2[6:0]) begin
          coeffs_65 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_66 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h42 == rs2[6:0]) begin
          coeffs_66 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_67 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h43 == rs2[6:0]) begin
          coeffs_67 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_68 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h44 == rs2[6:0]) begin
          coeffs_68 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_69 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h45 == rs2[6:0]) begin
          coeffs_69 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_70 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h46 == rs2[6:0]) begin
          coeffs_70 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_71 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h47 == rs2[6:0]) begin
          coeffs_71 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_72 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h48 == rs2[6:0]) begin
          coeffs_72 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_73 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h49 == rs2[6:0]) begin
          coeffs_73 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_74 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h4a == rs2[6:0]) begin
          coeffs_74 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_75 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h4b == rs2[6:0]) begin
          coeffs_75 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_76 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h4c == rs2[6:0]) begin
          coeffs_76 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_77 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h4d == rs2[6:0]) begin
          coeffs_77 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_78 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h4e == rs2[6:0]) begin
          coeffs_78 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_79 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h4f == rs2[6:0]) begin
          coeffs_79 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_80 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h50 == rs2[6:0]) begin
          coeffs_80 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_81 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h51 == rs2[6:0]) begin
          coeffs_81 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_82 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h52 == rs2[6:0]) begin
          coeffs_82 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_83 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h53 == rs2[6:0]) begin
          coeffs_83 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_84 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h54 == rs2[6:0]) begin
          coeffs_84 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_85 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h55 == rs2[6:0]) begin
          coeffs_85 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_86 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h56 == rs2[6:0]) begin
          coeffs_86 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_87 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h57 == rs2[6:0]) begin
          coeffs_87 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_88 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h58 == rs2[6:0]) begin
          coeffs_88 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_89 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h59 == rs2[6:0]) begin
          coeffs_89 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_90 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h5a == rs2[6:0]) begin
          coeffs_90 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_91 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h5b == rs2[6:0]) begin
          coeffs_91 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_92 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h5c == rs2[6:0]) begin
          coeffs_92 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_93 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h5d == rs2[6:0]) begin
          coeffs_93 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_94 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h5e == rs2[6:0]) begin
          coeffs_94 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_95 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h5f == rs2[6:0]) begin
          coeffs_95 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_96 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h60 == rs2[6:0]) begin
          coeffs_96 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_97 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h61 == rs2[6:0]) begin
          coeffs_97 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_98 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h62 == rs2[6:0]) begin
          coeffs_98 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_99 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (7'h63 == rs2[6:0]) begin
          coeffs_99 <= rs1;
        end
      end
    end
    if (reset) begin
      data_0 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_0 <= rs1;
        end
      end
    end
    if (reset) begin
      data_1 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_1 <= data_0;
        end
      end
    end
    if (reset) begin
      data_2 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_2 <= data_1;
        end
      end
    end
    if (reset) begin
      data_3 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_3 <= data_2;
        end
      end
    end
    if (reset) begin
      data_4 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_4 <= data_3;
        end
      end
    end
    if (reset) begin
      data_5 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_5 <= data_4;
        end
      end
    end
    if (reset) begin
      data_6 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_6 <= data_5;
        end
      end
    end
    if (reset) begin
      data_7 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_7 <= data_6;
        end
      end
    end
    if (reset) begin
      data_8 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_8 <= data_7;
        end
      end
    end
    if (reset) begin
      data_9 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_9 <= data_8;
        end
      end
    end
    if (reset) begin
      data_10 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_10 <= data_9;
        end
      end
    end
    if (reset) begin
      data_11 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_11 <= data_10;
        end
      end
    end
    if (reset) begin
      data_12 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_12 <= data_11;
        end
      end
    end
    if (reset) begin
      data_13 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_13 <= data_12;
        end
      end
    end
    if (reset) begin
      data_14 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_14 <= data_13;
        end
      end
    end
    if (reset) begin
      data_15 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_15 <= data_14;
        end
      end
    end
    if (reset) begin
      data_16 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_16 <= data_15;
        end
      end
    end
    if (reset) begin
      data_17 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_17 <= data_16;
        end
      end
    end
    if (reset) begin
      data_18 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_18 <= data_17;
        end
      end
    end
    if (reset) begin
      data_19 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_19 <= data_18;
        end
      end
    end
    if (reset) begin
      data_20 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_20 <= data_19;
        end
      end
    end
    if (reset) begin
      data_21 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_21 <= data_20;
        end
      end
    end
    if (reset) begin
      data_22 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_22 <= data_21;
        end
      end
    end
    if (reset) begin
      data_23 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_23 <= data_22;
        end
      end
    end
    if (reset) begin
      data_24 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_24 <= data_23;
        end
      end
    end
    if (reset) begin
      data_25 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_25 <= data_24;
        end
      end
    end
    if (reset) begin
      data_26 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_26 <= data_25;
        end
      end
    end
    if (reset) begin
      data_27 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_27 <= data_26;
        end
      end
    end
    if (reset) begin
      data_28 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_28 <= data_27;
        end
      end
    end
    if (reset) begin
      data_29 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_29 <= data_28;
        end
      end
    end
    if (reset) begin
      data_30 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_30 <= data_29;
        end
      end
    end
    if (reset) begin
      data_31 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_31 <= data_30;
        end
      end
    end
    if (reset) begin
      data_32 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_32 <= data_31;
        end
      end
    end
    if (reset) begin
      data_33 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_33 <= data_32;
        end
      end
    end
    if (reset) begin
      data_34 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_34 <= data_33;
        end
      end
    end
    if (reset) begin
      data_35 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_35 <= data_34;
        end
      end
    end
    if (reset) begin
      data_36 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_36 <= data_35;
        end
      end
    end
    if (reset) begin
      data_37 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_37 <= data_36;
        end
      end
    end
    if (reset) begin
      data_38 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_38 <= data_37;
        end
      end
    end
    if (reset) begin
      data_39 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_39 <= data_38;
        end
      end
    end
    if (reset) begin
      data_40 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_40 <= data_39;
        end
      end
    end
    if (reset) begin
      data_41 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_41 <= data_40;
        end
      end
    end
    if (reset) begin
      data_42 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_42 <= data_41;
        end
      end
    end
    if (reset) begin
      data_43 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_43 <= data_42;
        end
      end
    end
    if (reset) begin
      data_44 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_44 <= data_43;
        end
      end
    end
    if (reset) begin
      data_45 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_45 <= data_44;
        end
      end
    end
    if (reset) begin
      data_46 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_46 <= data_45;
        end
      end
    end
    if (reset) begin
      data_47 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_47 <= data_46;
        end
      end
    end
    if (reset) begin
      data_48 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_48 <= data_47;
        end
      end
    end
    if (reset) begin
      data_49 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_49 <= data_48;
        end
      end
    end
    if (reset) begin
      data_50 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_50 <= data_49;
        end
      end
    end
    if (reset) begin
      data_51 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_51 <= data_50;
        end
      end
    end
    if (reset) begin
      data_52 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_52 <= data_51;
        end
      end
    end
    if (reset) begin
      data_53 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_53 <= data_52;
        end
      end
    end
    if (reset) begin
      data_54 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_54 <= data_53;
        end
      end
    end
    if (reset) begin
      data_55 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_55 <= data_54;
        end
      end
    end
    if (reset) begin
      data_56 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_56 <= data_55;
        end
      end
    end
    if (reset) begin
      data_57 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_57 <= data_56;
        end
      end
    end
    if (reset) begin
      data_58 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_58 <= data_57;
        end
      end
    end
    if (reset) begin
      data_59 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_59 <= data_58;
        end
      end
    end
    if (reset) begin
      data_60 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_60 <= data_59;
        end
      end
    end
    if (reset) begin
      data_61 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_61 <= data_60;
        end
      end
    end
    if (reset) begin
      data_62 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_62 <= data_61;
        end
      end
    end
    if (reset) begin
      data_63 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_63 <= data_62;
        end
      end
    end
    if (reset) begin
      data_64 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_64 <= data_63;
        end
      end
    end
    if (reset) begin
      data_65 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_65 <= data_64;
        end
      end
    end
    if (reset) begin
      data_66 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_66 <= data_65;
        end
      end
    end
    if (reset) begin
      data_67 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_67 <= data_66;
        end
      end
    end
    if (reset) begin
      data_68 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_68 <= data_67;
        end
      end
    end
    if (reset) begin
      data_69 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_69 <= data_68;
        end
      end
    end
    if (reset) begin
      data_70 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_70 <= data_69;
        end
      end
    end
    if (reset) begin
      data_71 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_71 <= data_70;
        end
      end
    end
    if (reset) begin
      data_72 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_72 <= data_71;
        end
      end
    end
    if (reset) begin
      data_73 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_73 <= data_72;
        end
      end
    end
    if (reset) begin
      data_74 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_74 <= data_73;
        end
      end
    end
    if (reset) begin
      data_75 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_75 <= data_74;
        end
      end
    end
    if (reset) begin
      data_76 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_76 <= data_75;
        end
      end
    end
    if (reset) begin
      data_77 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_77 <= data_76;
        end
      end
    end
    if (reset) begin
      data_78 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_78 <= data_77;
        end
      end
    end
    if (reset) begin
      data_79 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_79 <= data_78;
        end
      end
    end
    if (reset) begin
      data_80 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_80 <= data_79;
        end
      end
    end
    if (reset) begin
      data_81 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_81 <= data_80;
        end
      end
    end
    if (reset) begin
      data_82 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_82 <= data_81;
        end
      end
    end
    if (reset) begin
      data_83 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_83 <= data_82;
        end
      end
    end
    if (reset) begin
      data_84 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_84 <= data_83;
        end
      end
    end
    if (reset) begin
      data_85 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_85 <= data_84;
        end
      end
    end
    if (reset) begin
      data_86 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_86 <= data_85;
        end
      end
    end
    if (reset) begin
      data_87 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_87 <= data_86;
        end
      end
    end
    if (reset) begin
      data_88 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_88 <= data_87;
        end
      end
    end
    if (reset) begin
      data_89 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_89 <= data_88;
        end
      end
    end
    if (reset) begin
      data_90 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_90 <= data_89;
        end
      end
    end
    if (reset) begin
      data_91 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_91 <= data_90;
        end
      end
    end
    if (reset) begin
      data_92 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_92 <= data_91;
        end
      end
    end
    if (reset) begin
      data_93 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_93 <= data_92;
        end
      end
    end
    if (reset) begin
      data_94 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_94 <= data_93;
        end
      end
    end
    if (reset) begin
      data_95 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_95 <= data_94;
        end
      end
    end
    if (reset) begin
      data_96 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_96 <= data_95;
        end
      end
    end
    if (reset) begin
      data_97 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_97 <= data_96;
        end
      end
    end
    if (reset) begin
      data_98 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_98 <= data_97;
        end
      end
    end
    if (reset) begin
      data_99 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_99 <= data_98;
        end
      end
    end
    if (reset) begin
      result <= 64'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        result <= {{32'd0}, _GEN_199};
      end else if (insn[6:0] == 7'h2b) begin
        result <= {{32'd0}, data_0};
      end else begin
        result <= _GEN_200;
      end
    end
  end
endmodule
