module SCIEPipelined #(parameter XLEN = 32)(
  input         clock,
  input         reset,
  input         valid,
  input  [31:0] insn,
  input  [31:0] rs1,
  input  [31:0] rs2,
  output [31:0] rd
);
  reg [31:0] coeffs_0;
  reg [31:0] coeffs_1;
  reg [31:0] coeffs_2;
  reg [31:0] coeffs_3;
  reg [31:0] coeffs_4;
  reg [31:0] coeffs_5;
  reg [31:0] coeffs_6;
  reg [31:0] coeffs_7;
  reg [31:0] coeffs_8;
  reg [31:0] coeffs_9;
  reg [31:0] data_0;
  reg [31:0] data_1;
  reg [31:0] data_2;
  reg [31:0] data_3;
  reg [31:0] data_4;
  reg [31:0] data_5;
  reg [31:0] data_6;
  reg [31:0] data_7;
  reg [31:0] data_8;
  reg [31:0] data_9;
  reg [63:0] result;
  wire [31:0] _GEN_11 = 4'h1 == rs2[3:0] ? coeffs_1 : coeffs_0;
  wire [31:0] _GEN_12 = 4'h2 == rs2[3:0] ? coeffs_2 : _GEN_11;
  wire [31:0] _GEN_13 = 4'h3 == rs2[3:0] ? coeffs_3 : _GEN_12;
  wire [31:0] _GEN_14 = 4'h4 == rs2[3:0] ? coeffs_4 : _GEN_13;
  wire [31:0] _GEN_15 = 4'h5 == rs2[3:0] ? coeffs_5 : _GEN_14;
  wire [31:0] _GEN_16 = 4'h6 == rs2[3:0] ? coeffs_6 : _GEN_15;
  wire [31:0] _GEN_17 = 4'h7 == rs2[3:0] ? coeffs_7 : _GEN_16;
  wire [31:0] _GEN_18 = 4'h8 == rs2[3:0] ? coeffs_8 : _GEN_17;
  wire [31:0] _GEN_19 = 4'h9 == rs2[3:0] ? coeffs_9 : _GEN_18;
  wire [63:0] _result_T_1 = data_0 * coeffs_0;
  wire [63:0] _result_T_2 = data_1 * coeffs_1;
  wire [63:0] _result_T_3 = data_2 * coeffs_2;
  wire [63:0] _result_T_4 = data_3 * coeffs_3;
  wire [63:0] _result_T_5 = data_4 * coeffs_4;
  wire [63:0] _result_T_6 = data_5 * coeffs_5;
  wire [63:0] _result_T_7 = data_6 * coeffs_6;
  wire [63:0] _result_T_8 = data_7 * coeffs_7;
  wire [63:0] _result_T_9 = data_8 * coeffs_8;
  wire [63:0] _result_T_10 = data_9 * coeffs_9;
  wire [63:0] _result_T_12 = _result_T_1 + _result_T_2;
  wire [63:0] _result_T_14 = _result_T_12 + _result_T_3;
  wire [63:0] _result_T_16 = _result_T_14 + _result_T_4;
  wire [63:0] _result_T_18 = _result_T_16 + _result_T_5;
  wire [63:0] _result_T_20 = _result_T_18 + _result_T_6;
  wire [63:0] _result_T_22 = _result_T_20 + _result_T_7;
  wire [63:0] _result_T_24 = _result_T_22 + _result_T_8;
  wire [63:0] _result_T_26 = _result_T_24 + _result_T_9;
  wire [63:0] _result_T_28 = _result_T_26 + _result_T_10;
  wire [63:0] _GEN_20 = insn[6:0] == 7'h3b ? _result_T_28 : result;
  assign rd = result[31:0];
  always @(posedge clock) begin
    if (reset) begin
      coeffs_0 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (4'h0 == rs2[3:0]) begin
          coeffs_0 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_1 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (4'h1 == rs2[3:0]) begin
          coeffs_1 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_2 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (4'h2 == rs2[3:0]) begin
          coeffs_2 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_3 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (4'h3 == rs2[3:0]) begin
          coeffs_3 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_4 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (4'h4 == rs2[3:0]) begin
          coeffs_4 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_5 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (4'h5 == rs2[3:0]) begin
          coeffs_5 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_6 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (4'h6 == rs2[3:0]) begin
          coeffs_6 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_7 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (4'h7 == rs2[3:0]) begin
          coeffs_7 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_8 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (4'h8 == rs2[3:0]) begin
          coeffs_8 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_9 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (4'h9 == rs2[3:0]) begin
          coeffs_9 <= rs1;
        end
      end
    end
    if (reset) begin
      data_0 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_0 <= rs1;
        end
      end
    end
    if (reset) begin
      data_1 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_1 <= data_0;
        end
      end
    end
    if (reset) begin
      data_2 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_2 <= data_1;
        end
      end
    end
    if (reset) begin
      data_3 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_3 <= data_2;
        end
      end
    end
    if (reset) begin
      data_4 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_4 <= data_3;
        end
      end
    end
    if (reset) begin
      data_5 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_5 <= data_4;
        end
      end
    end
    if (reset) begin
      data_6 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_6 <= data_5;
        end
      end
    end
    if (reset) begin
      data_7 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_7 <= data_6;
        end
      end
    end
    if (reset) begin
      data_8 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_8 <= data_7;
        end
      end
    end
    if (reset) begin
      data_9 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_9 <= data_8;
        end
      end
    end
    if (reset) begin
      result <= 64'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        result <= {{32'd0}, _GEN_19};
      end else if (insn[6:0] == 7'h2b) begin
        result <= {{32'd0}, data_0};
      end else begin
        result <= _GEN_20;
      end
    end
  end
endmodule
