module SCIEPipelined #(parameter XLEN = 32)(
  input         clock,
  input         reset,
  input         valid,
  input  [31:0] insn,
  input  [31:0] rs1,
  input  [31:0] rs2,
  output [31:0] rd
);
  reg [31:0] coeffs_0;
  reg [31:0] coeffs_1;
  reg [31:0] coeffs_2;
  reg [31:0] coeffs_3;
  reg [31:0] coeffs_4;
  reg [31:0] coeffs_5;
  reg [31:0] coeffs_6;
  reg [31:0] coeffs_7;
  reg [31:0] coeffs_8;
  reg [31:0] coeffs_9;
  reg [31:0] coeffs_10;
  reg [31:0] coeffs_11;
  reg [31:0] coeffs_12;
  reg [31:0] coeffs_13;
  reg [31:0] coeffs_14;
  reg [31:0] coeffs_15;
  reg [31:0] coeffs_16;
  reg [31:0] coeffs_17;
  reg [31:0] coeffs_18;
  reg [31:0] coeffs_19;
  reg [31:0] coeffs_20;
  reg [31:0] coeffs_21;
  reg [31:0] coeffs_22;
  reg [31:0] coeffs_23;
  reg [31:0] coeffs_24;
  reg [31:0] coeffs_25;
  reg [31:0] coeffs_26;
  reg [31:0] coeffs_27;
  reg [31:0] coeffs_28;
  reg [31:0] coeffs_29;
  reg [31:0] coeffs_30;
  reg [31:0] coeffs_31;
  reg [31:0] coeffs_32;
  reg [31:0] coeffs_33;
  reg [31:0] coeffs_34;
  reg [31:0] coeffs_35;
  reg [31:0] coeffs_36;
  reg [31:0] coeffs_37;
  reg [31:0] coeffs_38;
  reg [31:0] coeffs_39;
  reg [31:0] coeffs_40;
  reg [31:0] coeffs_41;
  reg [31:0] coeffs_42;
  reg [31:0] coeffs_43;
  reg [31:0] coeffs_44;
  reg [31:0] coeffs_45;
  reg [31:0] coeffs_46;
  reg [31:0] coeffs_47;
  reg [31:0] coeffs_48;
  reg [31:0] coeffs_49;
  reg [31:0] coeffs_50;
  reg [31:0] coeffs_51;
  reg [31:0] coeffs_52;
  reg [31:0] coeffs_53;
  reg [31:0] coeffs_54;
  reg [31:0] coeffs_55;
  reg [31:0] coeffs_56;
  reg [31:0] coeffs_57;
  reg [31:0] coeffs_58;
  reg [31:0] coeffs_59;
  reg [31:0] coeffs_60;
  reg [31:0] coeffs_61;
  reg [31:0] coeffs_62;
  reg [31:0] coeffs_63;
  reg [31:0] coeffs_64;
  reg [31:0] coeffs_65;
  reg [31:0] coeffs_66;
  reg [31:0] coeffs_67;
  reg [31:0] coeffs_68;
  reg [31:0] coeffs_69;
  reg [31:0] coeffs_70;
  reg [31:0] coeffs_71;
  reg [31:0] coeffs_72;
  reg [31:0] coeffs_73;
  reg [31:0] coeffs_74;
  reg [31:0] coeffs_75;
  reg [31:0] coeffs_76;
  reg [31:0] coeffs_77;
  reg [31:0] coeffs_78;
  reg [31:0] coeffs_79;
  reg [31:0] coeffs_80;
  reg [31:0] coeffs_81;
  reg [31:0] coeffs_82;
  reg [31:0] coeffs_83;
  reg [31:0] coeffs_84;
  reg [31:0] coeffs_85;
  reg [31:0] coeffs_86;
  reg [31:0] coeffs_87;
  reg [31:0] coeffs_88;
  reg [31:0] coeffs_89;
  reg [31:0] coeffs_90;
  reg [31:0] coeffs_91;
  reg [31:0] coeffs_92;
  reg [31:0] coeffs_93;
  reg [31:0] coeffs_94;
  reg [31:0] coeffs_95;
  reg [31:0] coeffs_96;
  reg [31:0] coeffs_97;
  reg [31:0] coeffs_98;
  reg [31:0] coeffs_99;
  reg [31:0] coeffs_100;
  reg [31:0] coeffs_101;
  reg [31:0] coeffs_102;
  reg [31:0] coeffs_103;
  reg [31:0] coeffs_104;
  reg [31:0] coeffs_105;
  reg [31:0] coeffs_106;
  reg [31:0] coeffs_107;
  reg [31:0] coeffs_108;
  reg [31:0] coeffs_109;
  reg [31:0] coeffs_110;
  reg [31:0] coeffs_111;
  reg [31:0] coeffs_112;
  reg [31:0] coeffs_113;
  reg [31:0] coeffs_114;
  reg [31:0] coeffs_115;
  reg [31:0] coeffs_116;
  reg [31:0] coeffs_117;
  reg [31:0] coeffs_118;
  reg [31:0] coeffs_119;
  reg [31:0] coeffs_120;
  reg [31:0] coeffs_121;
  reg [31:0] coeffs_122;
  reg [31:0] coeffs_123;
  reg [31:0] coeffs_124;
  reg [31:0] coeffs_125;
  reg [31:0] coeffs_126;
  reg [31:0] coeffs_127;
  reg [31:0] coeffs_128;
  reg [31:0] coeffs_129;
  reg [31:0] coeffs_130;
  reg [31:0] coeffs_131;
  reg [31:0] coeffs_132;
  reg [31:0] coeffs_133;
  reg [31:0] coeffs_134;
  reg [31:0] coeffs_135;
  reg [31:0] coeffs_136;
  reg [31:0] coeffs_137;
  reg [31:0] coeffs_138;
  reg [31:0] coeffs_139;
  reg [31:0] coeffs_140;
  reg [31:0] coeffs_141;
  reg [31:0] coeffs_142;
  reg [31:0] coeffs_143;
  reg [31:0] coeffs_144;
  reg [31:0] coeffs_145;
  reg [31:0] coeffs_146;
  reg [31:0] coeffs_147;
  reg [31:0] coeffs_148;
  reg [31:0] coeffs_149;
  reg [31:0] coeffs_150;
  reg [31:0] coeffs_151;
  reg [31:0] coeffs_152;
  reg [31:0] coeffs_153;
  reg [31:0] coeffs_154;
  reg [31:0] coeffs_155;
  reg [31:0] coeffs_156;
  reg [31:0] coeffs_157;
  reg [31:0] coeffs_158;
  reg [31:0] coeffs_159;
  reg [31:0] coeffs_160;
  reg [31:0] coeffs_161;
  reg [31:0] coeffs_162;
  reg [31:0] coeffs_163;
  reg [31:0] coeffs_164;
  reg [31:0] coeffs_165;
  reg [31:0] coeffs_166;
  reg [31:0] coeffs_167;
  reg [31:0] coeffs_168;
  reg [31:0] coeffs_169;
  reg [31:0] coeffs_170;
  reg [31:0] coeffs_171;
  reg [31:0] coeffs_172;
  reg [31:0] coeffs_173;
  reg [31:0] coeffs_174;
  reg [31:0] coeffs_175;
  reg [31:0] coeffs_176;
  reg [31:0] coeffs_177;
  reg [31:0] coeffs_178;
  reg [31:0] coeffs_179;
  reg [31:0] coeffs_180;
  reg [31:0] coeffs_181;
  reg [31:0] coeffs_182;
  reg [31:0] coeffs_183;
  reg [31:0] coeffs_184;
  reg [31:0] coeffs_185;
  reg [31:0] coeffs_186;
  reg [31:0] coeffs_187;
  reg [31:0] coeffs_188;
  reg [31:0] coeffs_189;
  reg [31:0] coeffs_190;
  reg [31:0] coeffs_191;
  reg [31:0] coeffs_192;
  reg [31:0] coeffs_193;
  reg [31:0] coeffs_194;
  reg [31:0] coeffs_195;
  reg [31:0] coeffs_196;
  reg [31:0] coeffs_197;
  reg [31:0] coeffs_198;
  reg [31:0] coeffs_199;
  reg [31:0] coeffs_200;
  reg [31:0] coeffs_201;
  reg [31:0] coeffs_202;
  reg [31:0] coeffs_203;
  reg [31:0] coeffs_204;
  reg [31:0] coeffs_205;
  reg [31:0] coeffs_206;
  reg [31:0] coeffs_207;
  reg [31:0] coeffs_208;
  reg [31:0] coeffs_209;
  reg [31:0] coeffs_210;
  reg [31:0] coeffs_211;
  reg [31:0] coeffs_212;
  reg [31:0] coeffs_213;
  reg [31:0] coeffs_214;
  reg [31:0] coeffs_215;
  reg [31:0] coeffs_216;
  reg [31:0] coeffs_217;
  reg [31:0] coeffs_218;
  reg [31:0] coeffs_219;
  reg [31:0] coeffs_220;
  reg [31:0] coeffs_221;
  reg [31:0] coeffs_222;
  reg [31:0] coeffs_223;
  reg [31:0] coeffs_224;
  reg [31:0] coeffs_225;
  reg [31:0] coeffs_226;
  reg [31:0] coeffs_227;
  reg [31:0] coeffs_228;
  reg [31:0] coeffs_229;
  reg [31:0] coeffs_230;
  reg [31:0] coeffs_231;
  reg [31:0] coeffs_232;
  reg [31:0] coeffs_233;
  reg [31:0] coeffs_234;
  reg [31:0] coeffs_235;
  reg [31:0] coeffs_236;
  reg [31:0] coeffs_237;
  reg [31:0] coeffs_238;
  reg [31:0] coeffs_239;
  reg [31:0] coeffs_240;
  reg [31:0] coeffs_241;
  reg [31:0] coeffs_242;
  reg [31:0] coeffs_243;
  reg [31:0] coeffs_244;
  reg [31:0] coeffs_245;
  reg [31:0] coeffs_246;
  reg [31:0] coeffs_247;
  reg [31:0] coeffs_248;
  reg [31:0] coeffs_249;
  reg [31:0] coeffs_250;
  reg [31:0] coeffs_251;
  reg [31:0] coeffs_252;
  reg [31:0] coeffs_253;
  reg [31:0] coeffs_254;
  reg [31:0] coeffs_255;
  reg [31:0] coeffs_256;
  reg [31:0] coeffs_257;
  reg [31:0] coeffs_258;
  reg [31:0] coeffs_259;
  reg [31:0] coeffs_260;
  reg [31:0] coeffs_261;
  reg [31:0] coeffs_262;
  reg [31:0] coeffs_263;
  reg [31:0] coeffs_264;
  reg [31:0] coeffs_265;
  reg [31:0] coeffs_266;
  reg [31:0] coeffs_267;
  reg [31:0] coeffs_268;
  reg [31:0] coeffs_269;
  reg [31:0] coeffs_270;
  reg [31:0] coeffs_271;
  reg [31:0] coeffs_272;
  reg [31:0] coeffs_273;
  reg [31:0] coeffs_274;
  reg [31:0] coeffs_275;
  reg [31:0] coeffs_276;
  reg [31:0] coeffs_277;
  reg [31:0] coeffs_278;
  reg [31:0] coeffs_279;
  reg [31:0] coeffs_280;
  reg [31:0] coeffs_281;
  reg [31:0] coeffs_282;
  reg [31:0] coeffs_283;
  reg [31:0] coeffs_284;
  reg [31:0] coeffs_285;
  reg [31:0] coeffs_286;
  reg [31:0] coeffs_287;
  reg [31:0] coeffs_288;
  reg [31:0] coeffs_289;
  reg [31:0] coeffs_290;
  reg [31:0] coeffs_291;
  reg [31:0] coeffs_292;
  reg [31:0] coeffs_293;
  reg [31:0] coeffs_294;
  reg [31:0] coeffs_295;
  reg [31:0] coeffs_296;
  reg [31:0] coeffs_297;
  reg [31:0] coeffs_298;
  reg [31:0] coeffs_299;
  reg [31:0] coeffs_300;
  reg [31:0] coeffs_301;
  reg [31:0] coeffs_302;
  reg [31:0] coeffs_303;
  reg [31:0] coeffs_304;
  reg [31:0] coeffs_305;
  reg [31:0] coeffs_306;
  reg [31:0] coeffs_307;
  reg [31:0] coeffs_308;
  reg [31:0] coeffs_309;
  reg [31:0] coeffs_310;
  reg [31:0] coeffs_311;
  reg [31:0] coeffs_312;
  reg [31:0] coeffs_313;
  reg [31:0] coeffs_314;
  reg [31:0] coeffs_315;
  reg [31:0] coeffs_316;
  reg [31:0] coeffs_317;
  reg [31:0] coeffs_318;
  reg [31:0] coeffs_319;
  reg [31:0] coeffs_320;
  reg [31:0] coeffs_321;
  reg [31:0] coeffs_322;
  reg [31:0] coeffs_323;
  reg [31:0] coeffs_324;
  reg [31:0] coeffs_325;
  reg [31:0] coeffs_326;
  reg [31:0] coeffs_327;
  reg [31:0] coeffs_328;
  reg [31:0] coeffs_329;
  reg [31:0] coeffs_330;
  reg [31:0] coeffs_331;
  reg [31:0] coeffs_332;
  reg [31:0] coeffs_333;
  reg [31:0] coeffs_334;
  reg [31:0] coeffs_335;
  reg [31:0] coeffs_336;
  reg [31:0] coeffs_337;
  reg [31:0] coeffs_338;
  reg [31:0] coeffs_339;
  reg [31:0] coeffs_340;
  reg [31:0] coeffs_341;
  reg [31:0] coeffs_342;
  reg [31:0] coeffs_343;
  reg [31:0] coeffs_344;
  reg [31:0] coeffs_345;
  reg [31:0] coeffs_346;
  reg [31:0] coeffs_347;
  reg [31:0] coeffs_348;
  reg [31:0] coeffs_349;
  reg [31:0] coeffs_350;
  reg [31:0] coeffs_351;
  reg [31:0] coeffs_352;
  reg [31:0] coeffs_353;
  reg [31:0] coeffs_354;
  reg [31:0] coeffs_355;
  reg [31:0] coeffs_356;
  reg [31:0] coeffs_357;
  reg [31:0] coeffs_358;
  reg [31:0] coeffs_359;
  reg [31:0] coeffs_360;
  reg [31:0] coeffs_361;
  reg [31:0] coeffs_362;
  reg [31:0] coeffs_363;
  reg [31:0] coeffs_364;
  reg [31:0] coeffs_365;
  reg [31:0] coeffs_366;
  reg [31:0] coeffs_367;
  reg [31:0] coeffs_368;
  reg [31:0] coeffs_369;
  reg [31:0] coeffs_370;
  reg [31:0] coeffs_371;
  reg [31:0] coeffs_372;
  reg [31:0] coeffs_373;
  reg [31:0] coeffs_374;
  reg [31:0] coeffs_375;
  reg [31:0] coeffs_376;
  reg [31:0] coeffs_377;
  reg [31:0] coeffs_378;
  reg [31:0] coeffs_379;
  reg [31:0] coeffs_380;
  reg [31:0] coeffs_381;
  reg [31:0] coeffs_382;
  reg [31:0] coeffs_383;
  reg [31:0] coeffs_384;
  reg [31:0] coeffs_385;
  reg [31:0] coeffs_386;
  reg [31:0] coeffs_387;
  reg [31:0] coeffs_388;
  reg [31:0] coeffs_389;
  reg [31:0] coeffs_390;
  reg [31:0] coeffs_391;
  reg [31:0] coeffs_392;
  reg [31:0] coeffs_393;
  reg [31:0] coeffs_394;
  reg [31:0] coeffs_395;
  reg [31:0] coeffs_396;
  reg [31:0] coeffs_397;
  reg [31:0] coeffs_398;
  reg [31:0] coeffs_399;
  reg [31:0] coeffs_400;
  reg [31:0] coeffs_401;
  reg [31:0] coeffs_402;
  reg [31:0] coeffs_403;
  reg [31:0] coeffs_404;
  reg [31:0] coeffs_405;
  reg [31:0] coeffs_406;
  reg [31:0] coeffs_407;
  reg [31:0] coeffs_408;
  reg [31:0] coeffs_409;
  reg [31:0] coeffs_410;
  reg [31:0] coeffs_411;
  reg [31:0] coeffs_412;
  reg [31:0] coeffs_413;
  reg [31:0] coeffs_414;
  reg [31:0] coeffs_415;
  reg [31:0] coeffs_416;
  reg [31:0] coeffs_417;
  reg [31:0] coeffs_418;
  reg [31:0] coeffs_419;
  reg [31:0] coeffs_420;
  reg [31:0] coeffs_421;
  reg [31:0] coeffs_422;
  reg [31:0] coeffs_423;
  reg [31:0] coeffs_424;
  reg [31:0] coeffs_425;
  reg [31:0] coeffs_426;
  reg [31:0] coeffs_427;
  reg [31:0] coeffs_428;
  reg [31:0] coeffs_429;
  reg [31:0] coeffs_430;
  reg [31:0] coeffs_431;
  reg [31:0] coeffs_432;
  reg [31:0] coeffs_433;
  reg [31:0] coeffs_434;
  reg [31:0] coeffs_435;
  reg [31:0] coeffs_436;
  reg [31:0] coeffs_437;
  reg [31:0] coeffs_438;
  reg [31:0] coeffs_439;
  reg [31:0] coeffs_440;
  reg [31:0] coeffs_441;
  reg [31:0] coeffs_442;
  reg [31:0] coeffs_443;
  reg [31:0] coeffs_444;
  reg [31:0] coeffs_445;
  reg [31:0] coeffs_446;
  reg [31:0] coeffs_447;
  reg [31:0] coeffs_448;
  reg [31:0] coeffs_449;
  reg [31:0] coeffs_450;
  reg [31:0] coeffs_451;
  reg [31:0] coeffs_452;
  reg [31:0] coeffs_453;
  reg [31:0] coeffs_454;
  reg [31:0] coeffs_455;
  reg [31:0] coeffs_456;
  reg [31:0] coeffs_457;
  reg [31:0] coeffs_458;
  reg [31:0] coeffs_459;
  reg [31:0] coeffs_460;
  reg [31:0] coeffs_461;
  reg [31:0] coeffs_462;
  reg [31:0] coeffs_463;
  reg [31:0] coeffs_464;
  reg [31:0] coeffs_465;
  reg [31:0] coeffs_466;
  reg [31:0] coeffs_467;
  reg [31:0] coeffs_468;
  reg [31:0] coeffs_469;
  reg [31:0] coeffs_470;
  reg [31:0] coeffs_471;
  reg [31:0] coeffs_472;
  reg [31:0] coeffs_473;
  reg [31:0] coeffs_474;
  reg [31:0] coeffs_475;
  reg [31:0] coeffs_476;
  reg [31:0] coeffs_477;
  reg [31:0] coeffs_478;
  reg [31:0] coeffs_479;
  reg [31:0] coeffs_480;
  reg [31:0] coeffs_481;
  reg [31:0] coeffs_482;
  reg [31:0] coeffs_483;
  reg [31:0] coeffs_484;
  reg [31:0] coeffs_485;
  reg [31:0] coeffs_486;
  reg [31:0] coeffs_487;
  reg [31:0] coeffs_488;
  reg [31:0] coeffs_489;
  reg [31:0] coeffs_490;
  reg [31:0] coeffs_491;
  reg [31:0] coeffs_492;
  reg [31:0] coeffs_493;
  reg [31:0] coeffs_494;
  reg [31:0] coeffs_495;
  reg [31:0] coeffs_496;
  reg [31:0] coeffs_497;
  reg [31:0] coeffs_498;
  reg [31:0] coeffs_499;
  reg [31:0] coeffs_500;
  reg [31:0] coeffs_501;
  reg [31:0] coeffs_502;
  reg [31:0] coeffs_503;
  reg [31:0] coeffs_504;
  reg [31:0] coeffs_505;
  reg [31:0] coeffs_506;
  reg [31:0] coeffs_507;
  reg [31:0] coeffs_508;
  reg [31:0] coeffs_509;
  reg [31:0] coeffs_510;
  reg [31:0] coeffs_511;
  reg [31:0] coeffs_512;
  reg [31:0] coeffs_513;
  reg [31:0] coeffs_514;
  reg [31:0] coeffs_515;
  reg [31:0] coeffs_516;
  reg [31:0] coeffs_517;
  reg [31:0] coeffs_518;
  reg [31:0] coeffs_519;
  reg [31:0] coeffs_520;
  reg [31:0] coeffs_521;
  reg [31:0] coeffs_522;
  reg [31:0] coeffs_523;
  reg [31:0] coeffs_524;
  reg [31:0] coeffs_525;
  reg [31:0] coeffs_526;
  reg [31:0] coeffs_527;
  reg [31:0] coeffs_528;
  reg [31:0] coeffs_529;
  reg [31:0] coeffs_530;
  reg [31:0] coeffs_531;
  reg [31:0] coeffs_532;
  reg [31:0] coeffs_533;
  reg [31:0] coeffs_534;
  reg [31:0] coeffs_535;
  reg [31:0] coeffs_536;
  reg [31:0] coeffs_537;
  reg [31:0] coeffs_538;
  reg [31:0] coeffs_539;
  reg [31:0] coeffs_540;
  reg [31:0] coeffs_541;
  reg [31:0] coeffs_542;
  reg [31:0] coeffs_543;
  reg [31:0] coeffs_544;
  reg [31:0] coeffs_545;
  reg [31:0] coeffs_546;
  reg [31:0] coeffs_547;
  reg [31:0] coeffs_548;
  reg [31:0] coeffs_549;
  reg [31:0] coeffs_550;
  reg [31:0] coeffs_551;
  reg [31:0] coeffs_552;
  reg [31:0] coeffs_553;
  reg [31:0] coeffs_554;
  reg [31:0] coeffs_555;
  reg [31:0] coeffs_556;
  reg [31:0] coeffs_557;
  reg [31:0] coeffs_558;
  reg [31:0] coeffs_559;
  reg [31:0] coeffs_560;
  reg [31:0] coeffs_561;
  reg [31:0] coeffs_562;
  reg [31:0] coeffs_563;
  reg [31:0] coeffs_564;
  reg [31:0] coeffs_565;
  reg [31:0] coeffs_566;
  reg [31:0] coeffs_567;
  reg [31:0] coeffs_568;
  reg [31:0] coeffs_569;
  reg [31:0] coeffs_570;
  reg [31:0] coeffs_571;
  reg [31:0] coeffs_572;
  reg [31:0] coeffs_573;
  reg [31:0] coeffs_574;
  reg [31:0] coeffs_575;
  reg [31:0] coeffs_576;
  reg [31:0] coeffs_577;
  reg [31:0] coeffs_578;
  reg [31:0] coeffs_579;
  reg [31:0] coeffs_580;
  reg [31:0] coeffs_581;
  reg [31:0] coeffs_582;
  reg [31:0] coeffs_583;
  reg [31:0] coeffs_584;
  reg [31:0] coeffs_585;
  reg [31:0] coeffs_586;
  reg [31:0] coeffs_587;
  reg [31:0] coeffs_588;
  reg [31:0] coeffs_589;
  reg [31:0] coeffs_590;
  reg [31:0] coeffs_591;
  reg [31:0] coeffs_592;
  reg [31:0] coeffs_593;
  reg [31:0] coeffs_594;
  reg [31:0] coeffs_595;
  reg [31:0] coeffs_596;
  reg [31:0] coeffs_597;
  reg [31:0] coeffs_598;
  reg [31:0] coeffs_599;
  reg [31:0] coeffs_600;
  reg [31:0] coeffs_601;
  reg [31:0] coeffs_602;
  reg [31:0] coeffs_603;
  reg [31:0] coeffs_604;
  reg [31:0] coeffs_605;
  reg [31:0] coeffs_606;
  reg [31:0] coeffs_607;
  reg [31:0] coeffs_608;
  reg [31:0] coeffs_609;
  reg [31:0] coeffs_610;
  reg [31:0] coeffs_611;
  reg [31:0] coeffs_612;
  reg [31:0] coeffs_613;
  reg [31:0] coeffs_614;
  reg [31:0] coeffs_615;
  reg [31:0] coeffs_616;
  reg [31:0] coeffs_617;
  reg [31:0] coeffs_618;
  reg [31:0] coeffs_619;
  reg [31:0] coeffs_620;
  reg [31:0] coeffs_621;
  reg [31:0] coeffs_622;
  reg [31:0] coeffs_623;
  reg [31:0] coeffs_624;
  reg [31:0] coeffs_625;
  reg [31:0] coeffs_626;
  reg [31:0] coeffs_627;
  reg [31:0] coeffs_628;
  reg [31:0] coeffs_629;
  reg [31:0] coeffs_630;
  reg [31:0] coeffs_631;
  reg [31:0] coeffs_632;
  reg [31:0] coeffs_633;
  reg [31:0] coeffs_634;
  reg [31:0] coeffs_635;
  reg [31:0] coeffs_636;
  reg [31:0] coeffs_637;
  reg [31:0] coeffs_638;
  reg [31:0] coeffs_639;
  reg [31:0] coeffs_640;
  reg [31:0] coeffs_641;
  reg [31:0] coeffs_642;
  reg [31:0] coeffs_643;
  reg [31:0] coeffs_644;
  reg [31:0] coeffs_645;
  reg [31:0] coeffs_646;
  reg [31:0] coeffs_647;
  reg [31:0] coeffs_648;
  reg [31:0] coeffs_649;
  reg [31:0] coeffs_650;
  reg [31:0] coeffs_651;
  reg [31:0] coeffs_652;
  reg [31:0] coeffs_653;
  reg [31:0] coeffs_654;
  reg [31:0] coeffs_655;
  reg [31:0] coeffs_656;
  reg [31:0] coeffs_657;
  reg [31:0] coeffs_658;
  reg [31:0] coeffs_659;
  reg [31:0] coeffs_660;
  reg [31:0] coeffs_661;
  reg [31:0] coeffs_662;
  reg [31:0] coeffs_663;
  reg [31:0] coeffs_664;
  reg [31:0] coeffs_665;
  reg [31:0] coeffs_666;
  reg [31:0] coeffs_667;
  reg [31:0] coeffs_668;
  reg [31:0] coeffs_669;
  reg [31:0] coeffs_670;
  reg [31:0] coeffs_671;
  reg [31:0] coeffs_672;
  reg [31:0] coeffs_673;
  reg [31:0] coeffs_674;
  reg [31:0] coeffs_675;
  reg [31:0] coeffs_676;
  reg [31:0] coeffs_677;
  reg [31:0] coeffs_678;
  reg [31:0] coeffs_679;
  reg [31:0] coeffs_680;
  reg [31:0] coeffs_681;
  reg [31:0] coeffs_682;
  reg [31:0] coeffs_683;
  reg [31:0] coeffs_684;
  reg [31:0] coeffs_685;
  reg [31:0] coeffs_686;
  reg [31:0] coeffs_687;
  reg [31:0] coeffs_688;
  reg [31:0] coeffs_689;
  reg [31:0] coeffs_690;
  reg [31:0] coeffs_691;
  reg [31:0] coeffs_692;
  reg [31:0] coeffs_693;
  reg [31:0] coeffs_694;
  reg [31:0] coeffs_695;
  reg [31:0] coeffs_696;
  reg [31:0] coeffs_697;
  reg [31:0] coeffs_698;
  reg [31:0] coeffs_699;
  reg [31:0] coeffs_700;
  reg [31:0] coeffs_701;
  reg [31:0] coeffs_702;
  reg [31:0] coeffs_703;
  reg [31:0] coeffs_704;
  reg [31:0] coeffs_705;
  reg [31:0] coeffs_706;
  reg [31:0] coeffs_707;
  reg [31:0] coeffs_708;
  reg [31:0] coeffs_709;
  reg [31:0] coeffs_710;
  reg [31:0] coeffs_711;
  reg [31:0] coeffs_712;
  reg [31:0] coeffs_713;
  reg [31:0] coeffs_714;
  reg [31:0] coeffs_715;
  reg [31:0] coeffs_716;
  reg [31:0] coeffs_717;
  reg [31:0] coeffs_718;
  reg [31:0] coeffs_719;
  reg [31:0] coeffs_720;
  reg [31:0] coeffs_721;
  reg [31:0] coeffs_722;
  reg [31:0] coeffs_723;
  reg [31:0] coeffs_724;
  reg [31:0] coeffs_725;
  reg [31:0] coeffs_726;
  reg [31:0] coeffs_727;
  reg [31:0] coeffs_728;
  reg [31:0] coeffs_729;
  reg [31:0] coeffs_730;
  reg [31:0] coeffs_731;
  reg [31:0] coeffs_732;
  reg [31:0] coeffs_733;
  reg [31:0] coeffs_734;
  reg [31:0] coeffs_735;
  reg [31:0] coeffs_736;
  reg [31:0] coeffs_737;
  reg [31:0] coeffs_738;
  reg [31:0] coeffs_739;
  reg [31:0] coeffs_740;
  reg [31:0] coeffs_741;
  reg [31:0] coeffs_742;
  reg [31:0] coeffs_743;
  reg [31:0] coeffs_744;
  reg [31:0] coeffs_745;
  reg [31:0] coeffs_746;
  reg [31:0] coeffs_747;
  reg [31:0] coeffs_748;
  reg [31:0] coeffs_749;
  reg [31:0] coeffs_750;
  reg [31:0] coeffs_751;
  reg [31:0] coeffs_752;
  reg [31:0] coeffs_753;
  reg [31:0] coeffs_754;
  reg [31:0] coeffs_755;
  reg [31:0] coeffs_756;
  reg [31:0] coeffs_757;
  reg [31:0] coeffs_758;
  reg [31:0] coeffs_759;
  reg [31:0] coeffs_760;
  reg [31:0] coeffs_761;
  reg [31:0] coeffs_762;
  reg [31:0] coeffs_763;
  reg [31:0] coeffs_764;
  reg [31:0] coeffs_765;
  reg [31:0] coeffs_766;
  reg [31:0] coeffs_767;
  reg [31:0] coeffs_768;
  reg [31:0] coeffs_769;
  reg [31:0] coeffs_770;
  reg [31:0] coeffs_771;
  reg [31:0] coeffs_772;
  reg [31:0] coeffs_773;
  reg [31:0] coeffs_774;
  reg [31:0] coeffs_775;
  reg [31:0] coeffs_776;
  reg [31:0] coeffs_777;
  reg [31:0] coeffs_778;
  reg [31:0] coeffs_779;
  reg [31:0] coeffs_780;
  reg [31:0] coeffs_781;
  reg [31:0] coeffs_782;
  reg [31:0] coeffs_783;
  reg [31:0] coeffs_784;
  reg [31:0] coeffs_785;
  reg [31:0] coeffs_786;
  reg [31:0] coeffs_787;
  reg [31:0] coeffs_788;
  reg [31:0] coeffs_789;
  reg [31:0] coeffs_790;
  reg [31:0] coeffs_791;
  reg [31:0] coeffs_792;
  reg [31:0] coeffs_793;
  reg [31:0] coeffs_794;
  reg [31:0] coeffs_795;
  reg [31:0] coeffs_796;
  reg [31:0] coeffs_797;
  reg [31:0] coeffs_798;
  reg [31:0] coeffs_799;
  reg [31:0] coeffs_800;
  reg [31:0] coeffs_801;
  reg [31:0] coeffs_802;
  reg [31:0] coeffs_803;
  reg [31:0] coeffs_804;
  reg [31:0] coeffs_805;
  reg [31:0] coeffs_806;
  reg [31:0] coeffs_807;
  reg [31:0] coeffs_808;
  reg [31:0] coeffs_809;
  reg [31:0] coeffs_810;
  reg [31:0] coeffs_811;
  reg [31:0] coeffs_812;
  reg [31:0] coeffs_813;
  reg [31:0] coeffs_814;
  reg [31:0] coeffs_815;
  reg [31:0] coeffs_816;
  reg [31:0] coeffs_817;
  reg [31:0] coeffs_818;
  reg [31:0] coeffs_819;
  reg [31:0] coeffs_820;
  reg [31:0] coeffs_821;
  reg [31:0] coeffs_822;
  reg [31:0] coeffs_823;
  reg [31:0] coeffs_824;
  reg [31:0] coeffs_825;
  reg [31:0] coeffs_826;
  reg [31:0] coeffs_827;
  reg [31:0] coeffs_828;
  reg [31:0] coeffs_829;
  reg [31:0] coeffs_830;
  reg [31:0] coeffs_831;
  reg [31:0] coeffs_832;
  reg [31:0] coeffs_833;
  reg [31:0] coeffs_834;
  reg [31:0] coeffs_835;
  reg [31:0] coeffs_836;
  reg [31:0] coeffs_837;
  reg [31:0] coeffs_838;
  reg [31:0] coeffs_839;
  reg [31:0] coeffs_840;
  reg [31:0] coeffs_841;
  reg [31:0] coeffs_842;
  reg [31:0] coeffs_843;
  reg [31:0] coeffs_844;
  reg [31:0] coeffs_845;
  reg [31:0] coeffs_846;
  reg [31:0] coeffs_847;
  reg [31:0] coeffs_848;
  reg [31:0] coeffs_849;
  reg [31:0] coeffs_850;
  reg [31:0] coeffs_851;
  reg [31:0] coeffs_852;
  reg [31:0] coeffs_853;
  reg [31:0] coeffs_854;
  reg [31:0] coeffs_855;
  reg [31:0] coeffs_856;
  reg [31:0] coeffs_857;
  reg [31:0] coeffs_858;
  reg [31:0] coeffs_859;
  reg [31:0] coeffs_860;
  reg [31:0] coeffs_861;
  reg [31:0] coeffs_862;
  reg [31:0] coeffs_863;
  reg [31:0] coeffs_864;
  reg [31:0] coeffs_865;
  reg [31:0] coeffs_866;
  reg [31:0] coeffs_867;
  reg [31:0] coeffs_868;
  reg [31:0] coeffs_869;
  reg [31:0] coeffs_870;
  reg [31:0] coeffs_871;
  reg [31:0] coeffs_872;
  reg [31:0] coeffs_873;
  reg [31:0] coeffs_874;
  reg [31:0] coeffs_875;
  reg [31:0] coeffs_876;
  reg [31:0] coeffs_877;
  reg [31:0] coeffs_878;
  reg [31:0] coeffs_879;
  reg [31:0] coeffs_880;
  reg [31:0] coeffs_881;
  reg [31:0] coeffs_882;
  reg [31:0] coeffs_883;
  reg [31:0] coeffs_884;
  reg [31:0] coeffs_885;
  reg [31:0] coeffs_886;
  reg [31:0] coeffs_887;
  reg [31:0] coeffs_888;
  reg [31:0] coeffs_889;
  reg [31:0] coeffs_890;
  reg [31:0] coeffs_891;
  reg [31:0] coeffs_892;
  reg [31:0] coeffs_893;
  reg [31:0] coeffs_894;
  reg [31:0] coeffs_895;
  reg [31:0] coeffs_896;
  reg [31:0] coeffs_897;
  reg [31:0] coeffs_898;
  reg [31:0] coeffs_899;
  reg [31:0] coeffs_900;
  reg [31:0] coeffs_901;
  reg [31:0] coeffs_902;
  reg [31:0] coeffs_903;
  reg [31:0] coeffs_904;
  reg [31:0] coeffs_905;
  reg [31:0] coeffs_906;
  reg [31:0] coeffs_907;
  reg [31:0] coeffs_908;
  reg [31:0] coeffs_909;
  reg [31:0] coeffs_910;
  reg [31:0] coeffs_911;
  reg [31:0] coeffs_912;
  reg [31:0] coeffs_913;
  reg [31:0] coeffs_914;
  reg [31:0] coeffs_915;
  reg [31:0] coeffs_916;
  reg [31:0] coeffs_917;
  reg [31:0] coeffs_918;
  reg [31:0] coeffs_919;
  reg [31:0] coeffs_920;
  reg [31:0] coeffs_921;
  reg [31:0] coeffs_922;
  reg [31:0] coeffs_923;
  reg [31:0] coeffs_924;
  reg [31:0] coeffs_925;
  reg [31:0] coeffs_926;
  reg [31:0] coeffs_927;
  reg [31:0] coeffs_928;
  reg [31:0] coeffs_929;
  reg [31:0] coeffs_930;
  reg [31:0] coeffs_931;
  reg [31:0] coeffs_932;
  reg [31:0] coeffs_933;
  reg [31:0] coeffs_934;
  reg [31:0] coeffs_935;
  reg [31:0] coeffs_936;
  reg [31:0] coeffs_937;
  reg [31:0] coeffs_938;
  reg [31:0] coeffs_939;
  reg [31:0] coeffs_940;
  reg [31:0] coeffs_941;
  reg [31:0] coeffs_942;
  reg [31:0] coeffs_943;
  reg [31:0] coeffs_944;
  reg [31:0] coeffs_945;
  reg [31:0] coeffs_946;
  reg [31:0] coeffs_947;
  reg [31:0] coeffs_948;
  reg [31:0] coeffs_949;
  reg [31:0] coeffs_950;
  reg [31:0] coeffs_951;
  reg [31:0] coeffs_952;
  reg [31:0] coeffs_953;
  reg [31:0] coeffs_954;
  reg [31:0] coeffs_955;
  reg [31:0] coeffs_956;
  reg [31:0] coeffs_957;
  reg [31:0] coeffs_958;
  reg [31:0] coeffs_959;
  reg [31:0] coeffs_960;
  reg [31:0] coeffs_961;
  reg [31:0] coeffs_962;
  reg [31:0] coeffs_963;
  reg [31:0] coeffs_964;
  reg [31:0] coeffs_965;
  reg [31:0] coeffs_966;
  reg [31:0] coeffs_967;
  reg [31:0] coeffs_968;
  reg [31:0] coeffs_969;
  reg [31:0] coeffs_970;
  reg [31:0] coeffs_971;
  reg [31:0] coeffs_972;
  reg [31:0] coeffs_973;
  reg [31:0] coeffs_974;
  reg [31:0] coeffs_975;
  reg [31:0] coeffs_976;
  reg [31:0] coeffs_977;
  reg [31:0] coeffs_978;
  reg [31:0] coeffs_979;
  reg [31:0] coeffs_980;
  reg [31:0] coeffs_981;
  reg [31:0] coeffs_982;
  reg [31:0] coeffs_983;
  reg [31:0] coeffs_984;
  reg [31:0] coeffs_985;
  reg [31:0] coeffs_986;
  reg [31:0] coeffs_987;
  reg [31:0] coeffs_988;
  reg [31:0] coeffs_989;
  reg [31:0] coeffs_990;
  reg [31:0] coeffs_991;
  reg [31:0] coeffs_992;
  reg [31:0] coeffs_993;
  reg [31:0] coeffs_994;
  reg [31:0] coeffs_995;
  reg [31:0] coeffs_996;
  reg [31:0] coeffs_997;
  reg [31:0] coeffs_998;
  reg [31:0] coeffs_999;
  reg [31:0] data_0;
  reg [31:0] data_1;
  reg [31:0] data_2;
  reg [31:0] data_3;
  reg [31:0] data_4;
  reg [31:0] data_5;
  reg [31:0] data_6;
  reg [31:0] data_7;
  reg [31:0] data_8;
  reg [31:0] data_9;
  reg [31:0] data_10;
  reg [31:0] data_11;
  reg [31:0] data_12;
  reg [31:0] data_13;
  reg [31:0] data_14;
  reg [31:0] data_15;
  reg [31:0] data_16;
  reg [31:0] data_17;
  reg [31:0] data_18;
  reg [31:0] data_19;
  reg [31:0] data_20;
  reg [31:0] data_21;
  reg [31:0] data_22;
  reg [31:0] data_23;
  reg [31:0] data_24;
  reg [31:0] data_25;
  reg [31:0] data_26;
  reg [31:0] data_27;
  reg [31:0] data_28;
  reg [31:0] data_29;
  reg [31:0] data_30;
  reg [31:0] data_31;
  reg [31:0] data_32;
  reg [31:0] data_33;
  reg [31:0] data_34;
  reg [31:0] data_35;
  reg [31:0] data_36;
  reg [31:0] data_37;
  reg [31:0] data_38;
  reg [31:0] data_39;
  reg [31:0] data_40;
  reg [31:0] data_41;
  reg [31:0] data_42;
  reg [31:0] data_43;
  reg [31:0] data_44;
  reg [31:0] data_45;
  reg [31:0] data_46;
  reg [31:0] data_47;
  reg [31:0] data_48;
  reg [31:0] data_49;
  reg [31:0] data_50;
  reg [31:0] data_51;
  reg [31:0] data_52;
  reg [31:0] data_53;
  reg [31:0] data_54;
  reg [31:0] data_55;
  reg [31:0] data_56;
  reg [31:0] data_57;
  reg [31:0] data_58;
  reg [31:0] data_59;
  reg [31:0] data_60;
  reg [31:0] data_61;
  reg [31:0] data_62;
  reg [31:0] data_63;
  reg [31:0] data_64;
  reg [31:0] data_65;
  reg [31:0] data_66;
  reg [31:0] data_67;
  reg [31:0] data_68;
  reg [31:0] data_69;
  reg [31:0] data_70;
  reg [31:0] data_71;
  reg [31:0] data_72;
  reg [31:0] data_73;
  reg [31:0] data_74;
  reg [31:0] data_75;
  reg [31:0] data_76;
  reg [31:0] data_77;
  reg [31:0] data_78;
  reg [31:0] data_79;
  reg [31:0] data_80;
  reg [31:0] data_81;
  reg [31:0] data_82;
  reg [31:0] data_83;
  reg [31:0] data_84;
  reg [31:0] data_85;
  reg [31:0] data_86;
  reg [31:0] data_87;
  reg [31:0] data_88;
  reg [31:0] data_89;
  reg [31:0] data_90;
  reg [31:0] data_91;
  reg [31:0] data_92;
  reg [31:0] data_93;
  reg [31:0] data_94;
  reg [31:0] data_95;
  reg [31:0] data_96;
  reg [31:0] data_97;
  reg [31:0] data_98;
  reg [31:0] data_99;
  reg [31:0] data_100;
  reg [31:0] data_101;
  reg [31:0] data_102;
  reg [31:0] data_103;
  reg [31:0] data_104;
  reg [31:0] data_105;
  reg [31:0] data_106;
  reg [31:0] data_107;
  reg [31:0] data_108;
  reg [31:0] data_109;
  reg [31:0] data_110;
  reg [31:0] data_111;
  reg [31:0] data_112;
  reg [31:0] data_113;
  reg [31:0] data_114;
  reg [31:0] data_115;
  reg [31:0] data_116;
  reg [31:0] data_117;
  reg [31:0] data_118;
  reg [31:0] data_119;
  reg [31:0] data_120;
  reg [31:0] data_121;
  reg [31:0] data_122;
  reg [31:0] data_123;
  reg [31:0] data_124;
  reg [31:0] data_125;
  reg [31:0] data_126;
  reg [31:0] data_127;
  reg [31:0] data_128;
  reg [31:0] data_129;
  reg [31:0] data_130;
  reg [31:0] data_131;
  reg [31:0] data_132;
  reg [31:0] data_133;
  reg [31:0] data_134;
  reg [31:0] data_135;
  reg [31:0] data_136;
  reg [31:0] data_137;
  reg [31:0] data_138;
  reg [31:0] data_139;
  reg [31:0] data_140;
  reg [31:0] data_141;
  reg [31:0] data_142;
  reg [31:0] data_143;
  reg [31:0] data_144;
  reg [31:0] data_145;
  reg [31:0] data_146;
  reg [31:0] data_147;
  reg [31:0] data_148;
  reg [31:0] data_149;
  reg [31:0] data_150;
  reg [31:0] data_151;
  reg [31:0] data_152;
  reg [31:0] data_153;
  reg [31:0] data_154;
  reg [31:0] data_155;
  reg [31:0] data_156;
  reg [31:0] data_157;
  reg [31:0] data_158;
  reg [31:0] data_159;
  reg [31:0] data_160;
  reg [31:0] data_161;
  reg [31:0] data_162;
  reg [31:0] data_163;
  reg [31:0] data_164;
  reg [31:0] data_165;
  reg [31:0] data_166;
  reg [31:0] data_167;
  reg [31:0] data_168;
  reg [31:0] data_169;
  reg [31:0] data_170;
  reg [31:0] data_171;
  reg [31:0] data_172;
  reg [31:0] data_173;
  reg [31:0] data_174;
  reg [31:0] data_175;
  reg [31:0] data_176;
  reg [31:0] data_177;
  reg [31:0] data_178;
  reg [31:0] data_179;
  reg [31:0] data_180;
  reg [31:0] data_181;
  reg [31:0] data_182;
  reg [31:0] data_183;
  reg [31:0] data_184;
  reg [31:0] data_185;
  reg [31:0] data_186;
  reg [31:0] data_187;
  reg [31:0] data_188;
  reg [31:0] data_189;
  reg [31:0] data_190;
  reg [31:0] data_191;
  reg [31:0] data_192;
  reg [31:0] data_193;
  reg [31:0] data_194;
  reg [31:0] data_195;
  reg [31:0] data_196;
  reg [31:0] data_197;
  reg [31:0] data_198;
  reg [31:0] data_199;
  reg [31:0] data_200;
  reg [31:0] data_201;
  reg [31:0] data_202;
  reg [31:0] data_203;
  reg [31:0] data_204;
  reg [31:0] data_205;
  reg [31:0] data_206;
  reg [31:0] data_207;
  reg [31:0] data_208;
  reg [31:0] data_209;
  reg [31:0] data_210;
  reg [31:0] data_211;
  reg [31:0] data_212;
  reg [31:0] data_213;
  reg [31:0] data_214;
  reg [31:0] data_215;
  reg [31:0] data_216;
  reg [31:0] data_217;
  reg [31:0] data_218;
  reg [31:0] data_219;
  reg [31:0] data_220;
  reg [31:0] data_221;
  reg [31:0] data_222;
  reg [31:0] data_223;
  reg [31:0] data_224;
  reg [31:0] data_225;
  reg [31:0] data_226;
  reg [31:0] data_227;
  reg [31:0] data_228;
  reg [31:0] data_229;
  reg [31:0] data_230;
  reg [31:0] data_231;
  reg [31:0] data_232;
  reg [31:0] data_233;
  reg [31:0] data_234;
  reg [31:0] data_235;
  reg [31:0] data_236;
  reg [31:0] data_237;
  reg [31:0] data_238;
  reg [31:0] data_239;
  reg [31:0] data_240;
  reg [31:0] data_241;
  reg [31:0] data_242;
  reg [31:0] data_243;
  reg [31:0] data_244;
  reg [31:0] data_245;
  reg [31:0] data_246;
  reg [31:0] data_247;
  reg [31:0] data_248;
  reg [31:0] data_249;
  reg [31:0] data_250;
  reg [31:0] data_251;
  reg [31:0] data_252;
  reg [31:0] data_253;
  reg [31:0] data_254;
  reg [31:0] data_255;
  reg [31:0] data_256;
  reg [31:0] data_257;
  reg [31:0] data_258;
  reg [31:0] data_259;
  reg [31:0] data_260;
  reg [31:0] data_261;
  reg [31:0] data_262;
  reg [31:0] data_263;
  reg [31:0] data_264;
  reg [31:0] data_265;
  reg [31:0] data_266;
  reg [31:0] data_267;
  reg [31:0] data_268;
  reg [31:0] data_269;
  reg [31:0] data_270;
  reg [31:0] data_271;
  reg [31:0] data_272;
  reg [31:0] data_273;
  reg [31:0] data_274;
  reg [31:0] data_275;
  reg [31:0] data_276;
  reg [31:0] data_277;
  reg [31:0] data_278;
  reg [31:0] data_279;
  reg [31:0] data_280;
  reg [31:0] data_281;
  reg [31:0] data_282;
  reg [31:0] data_283;
  reg [31:0] data_284;
  reg [31:0] data_285;
  reg [31:0] data_286;
  reg [31:0] data_287;
  reg [31:0] data_288;
  reg [31:0] data_289;
  reg [31:0] data_290;
  reg [31:0] data_291;
  reg [31:0] data_292;
  reg [31:0] data_293;
  reg [31:0] data_294;
  reg [31:0] data_295;
  reg [31:0] data_296;
  reg [31:0] data_297;
  reg [31:0] data_298;
  reg [31:0] data_299;
  reg [31:0] data_300;
  reg [31:0] data_301;
  reg [31:0] data_302;
  reg [31:0] data_303;
  reg [31:0] data_304;
  reg [31:0] data_305;
  reg [31:0] data_306;
  reg [31:0] data_307;
  reg [31:0] data_308;
  reg [31:0] data_309;
  reg [31:0] data_310;
  reg [31:0] data_311;
  reg [31:0] data_312;
  reg [31:0] data_313;
  reg [31:0] data_314;
  reg [31:0] data_315;
  reg [31:0] data_316;
  reg [31:0] data_317;
  reg [31:0] data_318;
  reg [31:0] data_319;
  reg [31:0] data_320;
  reg [31:0] data_321;
  reg [31:0] data_322;
  reg [31:0] data_323;
  reg [31:0] data_324;
  reg [31:0] data_325;
  reg [31:0] data_326;
  reg [31:0] data_327;
  reg [31:0] data_328;
  reg [31:0] data_329;
  reg [31:0] data_330;
  reg [31:0] data_331;
  reg [31:0] data_332;
  reg [31:0] data_333;
  reg [31:0] data_334;
  reg [31:0] data_335;
  reg [31:0] data_336;
  reg [31:0] data_337;
  reg [31:0] data_338;
  reg [31:0] data_339;
  reg [31:0] data_340;
  reg [31:0] data_341;
  reg [31:0] data_342;
  reg [31:0] data_343;
  reg [31:0] data_344;
  reg [31:0] data_345;
  reg [31:0] data_346;
  reg [31:0] data_347;
  reg [31:0] data_348;
  reg [31:0] data_349;
  reg [31:0] data_350;
  reg [31:0] data_351;
  reg [31:0] data_352;
  reg [31:0] data_353;
  reg [31:0] data_354;
  reg [31:0] data_355;
  reg [31:0] data_356;
  reg [31:0] data_357;
  reg [31:0] data_358;
  reg [31:0] data_359;
  reg [31:0] data_360;
  reg [31:0] data_361;
  reg [31:0] data_362;
  reg [31:0] data_363;
  reg [31:0] data_364;
  reg [31:0] data_365;
  reg [31:0] data_366;
  reg [31:0] data_367;
  reg [31:0] data_368;
  reg [31:0] data_369;
  reg [31:0] data_370;
  reg [31:0] data_371;
  reg [31:0] data_372;
  reg [31:0] data_373;
  reg [31:0] data_374;
  reg [31:0] data_375;
  reg [31:0] data_376;
  reg [31:0] data_377;
  reg [31:0] data_378;
  reg [31:0] data_379;
  reg [31:0] data_380;
  reg [31:0] data_381;
  reg [31:0] data_382;
  reg [31:0] data_383;
  reg [31:0] data_384;
  reg [31:0] data_385;
  reg [31:0] data_386;
  reg [31:0] data_387;
  reg [31:0] data_388;
  reg [31:0] data_389;
  reg [31:0] data_390;
  reg [31:0] data_391;
  reg [31:0] data_392;
  reg [31:0] data_393;
  reg [31:0] data_394;
  reg [31:0] data_395;
  reg [31:0] data_396;
  reg [31:0] data_397;
  reg [31:0] data_398;
  reg [31:0] data_399;
  reg [31:0] data_400;
  reg [31:0] data_401;
  reg [31:0] data_402;
  reg [31:0] data_403;
  reg [31:0] data_404;
  reg [31:0] data_405;
  reg [31:0] data_406;
  reg [31:0] data_407;
  reg [31:0] data_408;
  reg [31:0] data_409;
  reg [31:0] data_410;
  reg [31:0] data_411;
  reg [31:0] data_412;
  reg [31:0] data_413;
  reg [31:0] data_414;
  reg [31:0] data_415;
  reg [31:0] data_416;
  reg [31:0] data_417;
  reg [31:0] data_418;
  reg [31:0] data_419;
  reg [31:0] data_420;
  reg [31:0] data_421;
  reg [31:0] data_422;
  reg [31:0] data_423;
  reg [31:0] data_424;
  reg [31:0] data_425;
  reg [31:0] data_426;
  reg [31:0] data_427;
  reg [31:0] data_428;
  reg [31:0] data_429;
  reg [31:0] data_430;
  reg [31:0] data_431;
  reg [31:0] data_432;
  reg [31:0] data_433;
  reg [31:0] data_434;
  reg [31:0] data_435;
  reg [31:0] data_436;
  reg [31:0] data_437;
  reg [31:0] data_438;
  reg [31:0] data_439;
  reg [31:0] data_440;
  reg [31:0] data_441;
  reg [31:0] data_442;
  reg [31:0] data_443;
  reg [31:0] data_444;
  reg [31:0] data_445;
  reg [31:0] data_446;
  reg [31:0] data_447;
  reg [31:0] data_448;
  reg [31:0] data_449;
  reg [31:0] data_450;
  reg [31:0] data_451;
  reg [31:0] data_452;
  reg [31:0] data_453;
  reg [31:0] data_454;
  reg [31:0] data_455;
  reg [31:0] data_456;
  reg [31:0] data_457;
  reg [31:0] data_458;
  reg [31:0] data_459;
  reg [31:0] data_460;
  reg [31:0] data_461;
  reg [31:0] data_462;
  reg [31:0] data_463;
  reg [31:0] data_464;
  reg [31:0] data_465;
  reg [31:0] data_466;
  reg [31:0] data_467;
  reg [31:0] data_468;
  reg [31:0] data_469;
  reg [31:0] data_470;
  reg [31:0] data_471;
  reg [31:0] data_472;
  reg [31:0] data_473;
  reg [31:0] data_474;
  reg [31:0] data_475;
  reg [31:0] data_476;
  reg [31:0] data_477;
  reg [31:0] data_478;
  reg [31:0] data_479;
  reg [31:0] data_480;
  reg [31:0] data_481;
  reg [31:0] data_482;
  reg [31:0] data_483;
  reg [31:0] data_484;
  reg [31:0] data_485;
  reg [31:0] data_486;
  reg [31:0] data_487;
  reg [31:0] data_488;
  reg [31:0] data_489;
  reg [31:0] data_490;
  reg [31:0] data_491;
  reg [31:0] data_492;
  reg [31:0] data_493;
  reg [31:0] data_494;
  reg [31:0] data_495;
  reg [31:0] data_496;
  reg [31:0] data_497;
  reg [31:0] data_498;
  reg [31:0] data_499;
  reg [31:0] data_500;
  reg [31:0] data_501;
  reg [31:0] data_502;
  reg [31:0] data_503;
  reg [31:0] data_504;
  reg [31:0] data_505;
  reg [31:0] data_506;
  reg [31:0] data_507;
  reg [31:0] data_508;
  reg [31:0] data_509;
  reg [31:0] data_510;
  reg [31:0] data_511;
  reg [31:0] data_512;
  reg [31:0] data_513;
  reg [31:0] data_514;
  reg [31:0] data_515;
  reg [31:0] data_516;
  reg [31:0] data_517;
  reg [31:0] data_518;
  reg [31:0] data_519;
  reg [31:0] data_520;
  reg [31:0] data_521;
  reg [31:0] data_522;
  reg [31:0] data_523;
  reg [31:0] data_524;
  reg [31:0] data_525;
  reg [31:0] data_526;
  reg [31:0] data_527;
  reg [31:0] data_528;
  reg [31:0] data_529;
  reg [31:0] data_530;
  reg [31:0] data_531;
  reg [31:0] data_532;
  reg [31:0] data_533;
  reg [31:0] data_534;
  reg [31:0] data_535;
  reg [31:0] data_536;
  reg [31:0] data_537;
  reg [31:0] data_538;
  reg [31:0] data_539;
  reg [31:0] data_540;
  reg [31:0] data_541;
  reg [31:0] data_542;
  reg [31:0] data_543;
  reg [31:0] data_544;
  reg [31:0] data_545;
  reg [31:0] data_546;
  reg [31:0] data_547;
  reg [31:0] data_548;
  reg [31:0] data_549;
  reg [31:0] data_550;
  reg [31:0] data_551;
  reg [31:0] data_552;
  reg [31:0] data_553;
  reg [31:0] data_554;
  reg [31:0] data_555;
  reg [31:0] data_556;
  reg [31:0] data_557;
  reg [31:0] data_558;
  reg [31:0] data_559;
  reg [31:0] data_560;
  reg [31:0] data_561;
  reg [31:0] data_562;
  reg [31:0] data_563;
  reg [31:0] data_564;
  reg [31:0] data_565;
  reg [31:0] data_566;
  reg [31:0] data_567;
  reg [31:0] data_568;
  reg [31:0] data_569;
  reg [31:0] data_570;
  reg [31:0] data_571;
  reg [31:0] data_572;
  reg [31:0] data_573;
  reg [31:0] data_574;
  reg [31:0] data_575;
  reg [31:0] data_576;
  reg [31:0] data_577;
  reg [31:0] data_578;
  reg [31:0] data_579;
  reg [31:0] data_580;
  reg [31:0] data_581;
  reg [31:0] data_582;
  reg [31:0] data_583;
  reg [31:0] data_584;
  reg [31:0] data_585;
  reg [31:0] data_586;
  reg [31:0] data_587;
  reg [31:0] data_588;
  reg [31:0] data_589;
  reg [31:0] data_590;
  reg [31:0] data_591;
  reg [31:0] data_592;
  reg [31:0] data_593;
  reg [31:0] data_594;
  reg [31:0] data_595;
  reg [31:0] data_596;
  reg [31:0] data_597;
  reg [31:0] data_598;
  reg [31:0] data_599;
  reg [31:0] data_600;
  reg [31:0] data_601;
  reg [31:0] data_602;
  reg [31:0] data_603;
  reg [31:0] data_604;
  reg [31:0] data_605;
  reg [31:0] data_606;
  reg [31:0] data_607;
  reg [31:0] data_608;
  reg [31:0] data_609;
  reg [31:0] data_610;
  reg [31:0] data_611;
  reg [31:0] data_612;
  reg [31:0] data_613;
  reg [31:0] data_614;
  reg [31:0] data_615;
  reg [31:0] data_616;
  reg [31:0] data_617;
  reg [31:0] data_618;
  reg [31:0] data_619;
  reg [31:0] data_620;
  reg [31:0] data_621;
  reg [31:0] data_622;
  reg [31:0] data_623;
  reg [31:0] data_624;
  reg [31:0] data_625;
  reg [31:0] data_626;
  reg [31:0] data_627;
  reg [31:0] data_628;
  reg [31:0] data_629;
  reg [31:0] data_630;
  reg [31:0] data_631;
  reg [31:0] data_632;
  reg [31:0] data_633;
  reg [31:0] data_634;
  reg [31:0] data_635;
  reg [31:0] data_636;
  reg [31:0] data_637;
  reg [31:0] data_638;
  reg [31:0] data_639;
  reg [31:0] data_640;
  reg [31:0] data_641;
  reg [31:0] data_642;
  reg [31:0] data_643;
  reg [31:0] data_644;
  reg [31:0] data_645;
  reg [31:0] data_646;
  reg [31:0] data_647;
  reg [31:0] data_648;
  reg [31:0] data_649;
  reg [31:0] data_650;
  reg [31:0] data_651;
  reg [31:0] data_652;
  reg [31:0] data_653;
  reg [31:0] data_654;
  reg [31:0] data_655;
  reg [31:0] data_656;
  reg [31:0] data_657;
  reg [31:0] data_658;
  reg [31:0] data_659;
  reg [31:0] data_660;
  reg [31:0] data_661;
  reg [31:0] data_662;
  reg [31:0] data_663;
  reg [31:0] data_664;
  reg [31:0] data_665;
  reg [31:0] data_666;
  reg [31:0] data_667;
  reg [31:0] data_668;
  reg [31:0] data_669;
  reg [31:0] data_670;
  reg [31:0] data_671;
  reg [31:0] data_672;
  reg [31:0] data_673;
  reg [31:0] data_674;
  reg [31:0] data_675;
  reg [31:0] data_676;
  reg [31:0] data_677;
  reg [31:0] data_678;
  reg [31:0] data_679;
  reg [31:0] data_680;
  reg [31:0] data_681;
  reg [31:0] data_682;
  reg [31:0] data_683;
  reg [31:0] data_684;
  reg [31:0] data_685;
  reg [31:0] data_686;
  reg [31:0] data_687;
  reg [31:0] data_688;
  reg [31:0] data_689;
  reg [31:0] data_690;
  reg [31:0] data_691;
  reg [31:0] data_692;
  reg [31:0] data_693;
  reg [31:0] data_694;
  reg [31:0] data_695;
  reg [31:0] data_696;
  reg [31:0] data_697;
  reg [31:0] data_698;
  reg [31:0] data_699;
  reg [31:0] data_700;
  reg [31:0] data_701;
  reg [31:0] data_702;
  reg [31:0] data_703;
  reg [31:0] data_704;
  reg [31:0] data_705;
  reg [31:0] data_706;
  reg [31:0] data_707;
  reg [31:0] data_708;
  reg [31:0] data_709;
  reg [31:0] data_710;
  reg [31:0] data_711;
  reg [31:0] data_712;
  reg [31:0] data_713;
  reg [31:0] data_714;
  reg [31:0] data_715;
  reg [31:0] data_716;
  reg [31:0] data_717;
  reg [31:0] data_718;
  reg [31:0] data_719;
  reg [31:0] data_720;
  reg [31:0] data_721;
  reg [31:0] data_722;
  reg [31:0] data_723;
  reg [31:0] data_724;
  reg [31:0] data_725;
  reg [31:0] data_726;
  reg [31:0] data_727;
  reg [31:0] data_728;
  reg [31:0] data_729;
  reg [31:0] data_730;
  reg [31:0] data_731;
  reg [31:0] data_732;
  reg [31:0] data_733;
  reg [31:0] data_734;
  reg [31:0] data_735;
  reg [31:0] data_736;
  reg [31:0] data_737;
  reg [31:0] data_738;
  reg [31:0] data_739;
  reg [31:0] data_740;
  reg [31:0] data_741;
  reg [31:0] data_742;
  reg [31:0] data_743;
  reg [31:0] data_744;
  reg [31:0] data_745;
  reg [31:0] data_746;
  reg [31:0] data_747;
  reg [31:0] data_748;
  reg [31:0] data_749;
  reg [31:0] data_750;
  reg [31:0] data_751;
  reg [31:0] data_752;
  reg [31:0] data_753;
  reg [31:0] data_754;
  reg [31:0] data_755;
  reg [31:0] data_756;
  reg [31:0] data_757;
  reg [31:0] data_758;
  reg [31:0] data_759;
  reg [31:0] data_760;
  reg [31:0] data_761;
  reg [31:0] data_762;
  reg [31:0] data_763;
  reg [31:0] data_764;
  reg [31:0] data_765;
  reg [31:0] data_766;
  reg [31:0] data_767;
  reg [31:0] data_768;
  reg [31:0] data_769;
  reg [31:0] data_770;
  reg [31:0] data_771;
  reg [31:0] data_772;
  reg [31:0] data_773;
  reg [31:0] data_774;
  reg [31:0] data_775;
  reg [31:0] data_776;
  reg [31:0] data_777;
  reg [31:0] data_778;
  reg [31:0] data_779;
  reg [31:0] data_780;
  reg [31:0] data_781;
  reg [31:0] data_782;
  reg [31:0] data_783;
  reg [31:0] data_784;
  reg [31:0] data_785;
  reg [31:0] data_786;
  reg [31:0] data_787;
  reg [31:0] data_788;
  reg [31:0] data_789;
  reg [31:0] data_790;
  reg [31:0] data_791;
  reg [31:0] data_792;
  reg [31:0] data_793;
  reg [31:0] data_794;
  reg [31:0] data_795;
  reg [31:0] data_796;
  reg [31:0] data_797;
  reg [31:0] data_798;
  reg [31:0] data_799;
  reg [31:0] data_800;
  reg [31:0] data_801;
  reg [31:0] data_802;
  reg [31:0] data_803;
  reg [31:0] data_804;
  reg [31:0] data_805;
  reg [31:0] data_806;
  reg [31:0] data_807;
  reg [31:0] data_808;
  reg [31:0] data_809;
  reg [31:0] data_810;
  reg [31:0] data_811;
  reg [31:0] data_812;
  reg [31:0] data_813;
  reg [31:0] data_814;
  reg [31:0] data_815;
  reg [31:0] data_816;
  reg [31:0] data_817;
  reg [31:0] data_818;
  reg [31:0] data_819;
  reg [31:0] data_820;
  reg [31:0] data_821;
  reg [31:0] data_822;
  reg [31:0] data_823;
  reg [31:0] data_824;
  reg [31:0] data_825;
  reg [31:0] data_826;
  reg [31:0] data_827;
  reg [31:0] data_828;
  reg [31:0] data_829;
  reg [31:0] data_830;
  reg [31:0] data_831;
  reg [31:0] data_832;
  reg [31:0] data_833;
  reg [31:0] data_834;
  reg [31:0] data_835;
  reg [31:0] data_836;
  reg [31:0] data_837;
  reg [31:0] data_838;
  reg [31:0] data_839;
  reg [31:0] data_840;
  reg [31:0] data_841;
  reg [31:0] data_842;
  reg [31:0] data_843;
  reg [31:0] data_844;
  reg [31:0] data_845;
  reg [31:0] data_846;
  reg [31:0] data_847;
  reg [31:0] data_848;
  reg [31:0] data_849;
  reg [31:0] data_850;
  reg [31:0] data_851;
  reg [31:0] data_852;
  reg [31:0] data_853;
  reg [31:0] data_854;
  reg [31:0] data_855;
  reg [31:0] data_856;
  reg [31:0] data_857;
  reg [31:0] data_858;
  reg [31:0] data_859;
  reg [31:0] data_860;
  reg [31:0] data_861;
  reg [31:0] data_862;
  reg [31:0] data_863;
  reg [31:0] data_864;
  reg [31:0] data_865;
  reg [31:0] data_866;
  reg [31:0] data_867;
  reg [31:0] data_868;
  reg [31:0] data_869;
  reg [31:0] data_870;
  reg [31:0] data_871;
  reg [31:0] data_872;
  reg [31:0] data_873;
  reg [31:0] data_874;
  reg [31:0] data_875;
  reg [31:0] data_876;
  reg [31:0] data_877;
  reg [31:0] data_878;
  reg [31:0] data_879;
  reg [31:0] data_880;
  reg [31:0] data_881;
  reg [31:0] data_882;
  reg [31:0] data_883;
  reg [31:0] data_884;
  reg [31:0] data_885;
  reg [31:0] data_886;
  reg [31:0] data_887;
  reg [31:0] data_888;
  reg [31:0] data_889;
  reg [31:0] data_890;
  reg [31:0] data_891;
  reg [31:0] data_892;
  reg [31:0] data_893;
  reg [31:0] data_894;
  reg [31:0] data_895;
  reg [31:0] data_896;
  reg [31:0] data_897;
  reg [31:0] data_898;
  reg [31:0] data_899;
  reg [31:0] data_900;
  reg [31:0] data_901;
  reg [31:0] data_902;
  reg [31:0] data_903;
  reg [31:0] data_904;
  reg [31:0] data_905;
  reg [31:0] data_906;
  reg [31:0] data_907;
  reg [31:0] data_908;
  reg [31:0] data_909;
  reg [31:0] data_910;
  reg [31:0] data_911;
  reg [31:0] data_912;
  reg [31:0] data_913;
  reg [31:0] data_914;
  reg [31:0] data_915;
  reg [31:0] data_916;
  reg [31:0] data_917;
  reg [31:0] data_918;
  reg [31:0] data_919;
  reg [31:0] data_920;
  reg [31:0] data_921;
  reg [31:0] data_922;
  reg [31:0] data_923;
  reg [31:0] data_924;
  reg [31:0] data_925;
  reg [31:0] data_926;
  reg [31:0] data_927;
  reg [31:0] data_928;
  reg [31:0] data_929;
  reg [31:0] data_930;
  reg [31:0] data_931;
  reg [31:0] data_932;
  reg [31:0] data_933;
  reg [31:0] data_934;
  reg [31:0] data_935;
  reg [31:0] data_936;
  reg [31:0] data_937;
  reg [31:0] data_938;
  reg [31:0] data_939;
  reg [31:0] data_940;
  reg [31:0] data_941;
  reg [31:0] data_942;
  reg [31:0] data_943;
  reg [31:0] data_944;
  reg [31:0] data_945;
  reg [31:0] data_946;
  reg [31:0] data_947;
  reg [31:0] data_948;
  reg [31:0] data_949;
  reg [31:0] data_950;
  reg [31:0] data_951;
  reg [31:0] data_952;
  reg [31:0] data_953;
  reg [31:0] data_954;
  reg [31:0] data_955;
  reg [31:0] data_956;
  reg [31:0] data_957;
  reg [31:0] data_958;
  reg [31:0] data_959;
  reg [31:0] data_960;
  reg [31:0] data_961;
  reg [31:0] data_962;
  reg [31:0] data_963;
  reg [31:0] data_964;
  reg [31:0] data_965;
  reg [31:0] data_966;
  reg [31:0] data_967;
  reg [31:0] data_968;
  reg [31:0] data_969;
  reg [31:0] data_970;
  reg [31:0] data_971;
  reg [31:0] data_972;
  reg [31:0] data_973;
  reg [31:0] data_974;
  reg [31:0] data_975;
  reg [31:0] data_976;
  reg [31:0] data_977;
  reg [31:0] data_978;
  reg [31:0] data_979;
  reg [31:0] data_980;
  reg [31:0] data_981;
  reg [31:0] data_982;
  reg [31:0] data_983;
  reg [31:0] data_984;
  reg [31:0] data_985;
  reg [31:0] data_986;
  reg [31:0] data_987;
  reg [31:0] data_988;
  reg [31:0] data_989;
  reg [31:0] data_990;
  reg [31:0] data_991;
  reg [31:0] data_992;
  reg [31:0] data_993;
  reg [31:0] data_994;
  reg [31:0] data_995;
  reg [31:0] data_996;
  reg [31:0] data_997;
  reg [31:0] data_998;
  reg [31:0] data_999;
  reg [63:0] result;
  wire [31:0] _GEN_1001 = 10'h1 == rs2[9:0] ? coeffs_1 : coeffs_0;
  wire [31:0] _GEN_1002 = 10'h2 == rs2[9:0] ? coeffs_2 : _GEN_1001;
  wire [31:0] _GEN_1003 = 10'h3 == rs2[9:0] ? coeffs_3 : _GEN_1002;
  wire [31:0] _GEN_1004 = 10'h4 == rs2[9:0] ? coeffs_4 : _GEN_1003;
  wire [31:0] _GEN_1005 = 10'h5 == rs2[9:0] ? coeffs_5 : _GEN_1004;
  wire [31:0] _GEN_1006 = 10'h6 == rs2[9:0] ? coeffs_6 : _GEN_1005;
  wire [31:0] _GEN_1007 = 10'h7 == rs2[9:0] ? coeffs_7 : _GEN_1006;
  wire [31:0] _GEN_1008 = 10'h8 == rs2[9:0] ? coeffs_8 : _GEN_1007;
  wire [31:0] _GEN_1009 = 10'h9 == rs2[9:0] ? coeffs_9 : _GEN_1008;
  wire [31:0] _GEN_1010 = 10'ha == rs2[9:0] ? coeffs_10 : _GEN_1009;
  wire [31:0] _GEN_1011 = 10'hb == rs2[9:0] ? coeffs_11 : _GEN_1010;
  wire [31:0] _GEN_1012 = 10'hc == rs2[9:0] ? coeffs_12 : _GEN_1011;
  wire [31:0] _GEN_1013 = 10'hd == rs2[9:0] ? coeffs_13 : _GEN_1012;
  wire [31:0] _GEN_1014 = 10'he == rs2[9:0] ? coeffs_14 : _GEN_1013;
  wire [31:0] _GEN_1015 = 10'hf == rs2[9:0] ? coeffs_15 : _GEN_1014;
  wire [31:0] _GEN_1016 = 10'h10 == rs2[9:0] ? coeffs_16 : _GEN_1015;
  wire [31:0] _GEN_1017 = 10'h11 == rs2[9:0] ? coeffs_17 : _GEN_1016;
  wire [31:0] _GEN_1018 = 10'h12 == rs2[9:0] ? coeffs_18 : _GEN_1017;
  wire [31:0] _GEN_1019 = 10'h13 == rs2[9:0] ? coeffs_19 : _GEN_1018;
  wire [31:0] _GEN_1020 = 10'h14 == rs2[9:0] ? coeffs_20 : _GEN_1019;
  wire [31:0] _GEN_1021 = 10'h15 == rs2[9:0] ? coeffs_21 : _GEN_1020;
  wire [31:0] _GEN_1022 = 10'h16 == rs2[9:0] ? coeffs_22 : _GEN_1021;
  wire [31:0] _GEN_1023 = 10'h17 == rs2[9:0] ? coeffs_23 : _GEN_1022;
  wire [31:0] _GEN_1024 = 10'h18 == rs2[9:0] ? coeffs_24 : _GEN_1023;
  wire [31:0] _GEN_1025 = 10'h19 == rs2[9:0] ? coeffs_25 : _GEN_1024;
  wire [31:0] _GEN_1026 = 10'h1a == rs2[9:0] ? coeffs_26 : _GEN_1025;
  wire [31:0] _GEN_1027 = 10'h1b == rs2[9:0] ? coeffs_27 : _GEN_1026;
  wire [31:0] _GEN_1028 = 10'h1c == rs2[9:0] ? coeffs_28 : _GEN_1027;
  wire [31:0] _GEN_1029 = 10'h1d == rs2[9:0] ? coeffs_29 : _GEN_1028;
  wire [31:0] _GEN_1030 = 10'h1e == rs2[9:0] ? coeffs_30 : _GEN_1029;
  wire [31:0] _GEN_1031 = 10'h1f == rs2[9:0] ? coeffs_31 : _GEN_1030;
  wire [31:0] _GEN_1032 = 10'h20 == rs2[9:0] ? coeffs_32 : _GEN_1031;
  wire [31:0] _GEN_1033 = 10'h21 == rs2[9:0] ? coeffs_33 : _GEN_1032;
  wire [31:0] _GEN_1034 = 10'h22 == rs2[9:0] ? coeffs_34 : _GEN_1033;
  wire [31:0] _GEN_1035 = 10'h23 == rs2[9:0] ? coeffs_35 : _GEN_1034;
  wire [31:0] _GEN_1036 = 10'h24 == rs2[9:0] ? coeffs_36 : _GEN_1035;
  wire [31:0] _GEN_1037 = 10'h25 == rs2[9:0] ? coeffs_37 : _GEN_1036;
  wire [31:0] _GEN_1038 = 10'h26 == rs2[9:0] ? coeffs_38 : _GEN_1037;
  wire [31:0] _GEN_1039 = 10'h27 == rs2[9:0] ? coeffs_39 : _GEN_1038;
  wire [31:0] _GEN_1040 = 10'h28 == rs2[9:0] ? coeffs_40 : _GEN_1039;
  wire [31:0] _GEN_1041 = 10'h29 == rs2[9:0] ? coeffs_41 : _GEN_1040;
  wire [31:0] _GEN_1042 = 10'h2a == rs2[9:0] ? coeffs_42 : _GEN_1041;
  wire [31:0] _GEN_1043 = 10'h2b == rs2[9:0] ? coeffs_43 : _GEN_1042;
  wire [31:0] _GEN_1044 = 10'h2c == rs2[9:0] ? coeffs_44 : _GEN_1043;
  wire [31:0] _GEN_1045 = 10'h2d == rs2[9:0] ? coeffs_45 : _GEN_1044;
  wire [31:0] _GEN_1046 = 10'h2e == rs2[9:0] ? coeffs_46 : _GEN_1045;
  wire [31:0] _GEN_1047 = 10'h2f == rs2[9:0] ? coeffs_47 : _GEN_1046;
  wire [31:0] _GEN_1048 = 10'h30 == rs2[9:0] ? coeffs_48 : _GEN_1047;
  wire [31:0] _GEN_1049 = 10'h31 == rs2[9:0] ? coeffs_49 : _GEN_1048;
  wire [31:0] _GEN_1050 = 10'h32 == rs2[9:0] ? coeffs_50 : _GEN_1049;
  wire [31:0] _GEN_1051 = 10'h33 == rs2[9:0] ? coeffs_51 : _GEN_1050;
  wire [31:0] _GEN_1052 = 10'h34 == rs2[9:0] ? coeffs_52 : _GEN_1051;
  wire [31:0] _GEN_1053 = 10'h35 == rs2[9:0] ? coeffs_53 : _GEN_1052;
  wire [31:0] _GEN_1054 = 10'h36 == rs2[9:0] ? coeffs_54 : _GEN_1053;
  wire [31:0] _GEN_1055 = 10'h37 == rs2[9:0] ? coeffs_55 : _GEN_1054;
  wire [31:0] _GEN_1056 = 10'h38 == rs2[9:0] ? coeffs_56 : _GEN_1055;
  wire [31:0] _GEN_1057 = 10'h39 == rs2[9:0] ? coeffs_57 : _GEN_1056;
  wire [31:0] _GEN_1058 = 10'h3a == rs2[9:0] ? coeffs_58 : _GEN_1057;
  wire [31:0] _GEN_1059 = 10'h3b == rs2[9:0] ? coeffs_59 : _GEN_1058;
  wire [31:0] _GEN_1060 = 10'h3c == rs2[9:0] ? coeffs_60 : _GEN_1059;
  wire [31:0] _GEN_1061 = 10'h3d == rs2[9:0] ? coeffs_61 : _GEN_1060;
  wire [31:0] _GEN_1062 = 10'h3e == rs2[9:0] ? coeffs_62 : _GEN_1061;
  wire [31:0] _GEN_1063 = 10'h3f == rs2[9:0] ? coeffs_63 : _GEN_1062;
  wire [31:0] _GEN_1064 = 10'h40 == rs2[9:0] ? coeffs_64 : _GEN_1063;
  wire [31:0] _GEN_1065 = 10'h41 == rs2[9:0] ? coeffs_65 : _GEN_1064;
  wire [31:0] _GEN_1066 = 10'h42 == rs2[9:0] ? coeffs_66 : _GEN_1065;
  wire [31:0] _GEN_1067 = 10'h43 == rs2[9:0] ? coeffs_67 : _GEN_1066;
  wire [31:0] _GEN_1068 = 10'h44 == rs2[9:0] ? coeffs_68 : _GEN_1067;
  wire [31:0] _GEN_1069 = 10'h45 == rs2[9:0] ? coeffs_69 : _GEN_1068;
  wire [31:0] _GEN_1070 = 10'h46 == rs2[9:0] ? coeffs_70 : _GEN_1069;
  wire [31:0] _GEN_1071 = 10'h47 == rs2[9:0] ? coeffs_71 : _GEN_1070;
  wire [31:0] _GEN_1072 = 10'h48 == rs2[9:0] ? coeffs_72 : _GEN_1071;
  wire [31:0] _GEN_1073 = 10'h49 == rs2[9:0] ? coeffs_73 : _GEN_1072;
  wire [31:0] _GEN_1074 = 10'h4a == rs2[9:0] ? coeffs_74 : _GEN_1073;
  wire [31:0] _GEN_1075 = 10'h4b == rs2[9:0] ? coeffs_75 : _GEN_1074;
  wire [31:0] _GEN_1076 = 10'h4c == rs2[9:0] ? coeffs_76 : _GEN_1075;
  wire [31:0] _GEN_1077 = 10'h4d == rs2[9:0] ? coeffs_77 : _GEN_1076;
  wire [31:0] _GEN_1078 = 10'h4e == rs2[9:0] ? coeffs_78 : _GEN_1077;
  wire [31:0] _GEN_1079 = 10'h4f == rs2[9:0] ? coeffs_79 : _GEN_1078;
  wire [31:0] _GEN_1080 = 10'h50 == rs2[9:0] ? coeffs_80 : _GEN_1079;
  wire [31:0] _GEN_1081 = 10'h51 == rs2[9:0] ? coeffs_81 : _GEN_1080;
  wire [31:0] _GEN_1082 = 10'h52 == rs2[9:0] ? coeffs_82 : _GEN_1081;
  wire [31:0] _GEN_1083 = 10'h53 == rs2[9:0] ? coeffs_83 : _GEN_1082;
  wire [31:0] _GEN_1084 = 10'h54 == rs2[9:0] ? coeffs_84 : _GEN_1083;
  wire [31:0] _GEN_1085 = 10'h55 == rs2[9:0] ? coeffs_85 : _GEN_1084;
  wire [31:0] _GEN_1086 = 10'h56 == rs2[9:0] ? coeffs_86 : _GEN_1085;
  wire [31:0] _GEN_1087 = 10'h57 == rs2[9:0] ? coeffs_87 : _GEN_1086;
  wire [31:0] _GEN_1088 = 10'h58 == rs2[9:0] ? coeffs_88 : _GEN_1087;
  wire [31:0] _GEN_1089 = 10'h59 == rs2[9:0] ? coeffs_89 : _GEN_1088;
  wire [31:0] _GEN_1090 = 10'h5a == rs2[9:0] ? coeffs_90 : _GEN_1089;
  wire [31:0] _GEN_1091 = 10'h5b == rs2[9:0] ? coeffs_91 : _GEN_1090;
  wire [31:0] _GEN_1092 = 10'h5c == rs2[9:0] ? coeffs_92 : _GEN_1091;
  wire [31:0] _GEN_1093 = 10'h5d == rs2[9:0] ? coeffs_93 : _GEN_1092;
  wire [31:0] _GEN_1094 = 10'h5e == rs2[9:0] ? coeffs_94 : _GEN_1093;
  wire [31:0] _GEN_1095 = 10'h5f == rs2[9:0] ? coeffs_95 : _GEN_1094;
  wire [31:0] _GEN_1096 = 10'h60 == rs2[9:0] ? coeffs_96 : _GEN_1095;
  wire [31:0] _GEN_1097 = 10'h61 == rs2[9:0] ? coeffs_97 : _GEN_1096;
  wire [31:0] _GEN_1098 = 10'h62 == rs2[9:0] ? coeffs_98 : _GEN_1097;
  wire [31:0] _GEN_1099 = 10'h63 == rs2[9:0] ? coeffs_99 : _GEN_1098;
  wire [31:0] _GEN_1100 = 10'h64 == rs2[9:0] ? coeffs_100 : _GEN_1099;
  wire [31:0] _GEN_1101 = 10'h65 == rs2[9:0] ? coeffs_101 : _GEN_1100;
  wire [31:0] _GEN_1102 = 10'h66 == rs2[9:0] ? coeffs_102 : _GEN_1101;
  wire [31:0] _GEN_1103 = 10'h67 == rs2[9:0] ? coeffs_103 : _GEN_1102;
  wire [31:0] _GEN_1104 = 10'h68 == rs2[9:0] ? coeffs_104 : _GEN_1103;
  wire [31:0] _GEN_1105 = 10'h69 == rs2[9:0] ? coeffs_105 : _GEN_1104;
  wire [31:0] _GEN_1106 = 10'h6a == rs2[9:0] ? coeffs_106 : _GEN_1105;
  wire [31:0] _GEN_1107 = 10'h6b == rs2[9:0] ? coeffs_107 : _GEN_1106;
  wire [31:0] _GEN_1108 = 10'h6c == rs2[9:0] ? coeffs_108 : _GEN_1107;
  wire [31:0] _GEN_1109 = 10'h6d == rs2[9:0] ? coeffs_109 : _GEN_1108;
  wire [31:0] _GEN_1110 = 10'h6e == rs2[9:0] ? coeffs_110 : _GEN_1109;
  wire [31:0] _GEN_1111 = 10'h6f == rs2[9:0] ? coeffs_111 : _GEN_1110;
  wire [31:0] _GEN_1112 = 10'h70 == rs2[9:0] ? coeffs_112 : _GEN_1111;
  wire [31:0] _GEN_1113 = 10'h71 == rs2[9:0] ? coeffs_113 : _GEN_1112;
  wire [31:0] _GEN_1114 = 10'h72 == rs2[9:0] ? coeffs_114 : _GEN_1113;
  wire [31:0] _GEN_1115 = 10'h73 == rs2[9:0] ? coeffs_115 : _GEN_1114;
  wire [31:0] _GEN_1116 = 10'h74 == rs2[9:0] ? coeffs_116 : _GEN_1115;
  wire [31:0] _GEN_1117 = 10'h75 == rs2[9:0] ? coeffs_117 : _GEN_1116;
  wire [31:0] _GEN_1118 = 10'h76 == rs2[9:0] ? coeffs_118 : _GEN_1117;
  wire [31:0] _GEN_1119 = 10'h77 == rs2[9:0] ? coeffs_119 : _GEN_1118;
  wire [31:0] _GEN_1120 = 10'h78 == rs2[9:0] ? coeffs_120 : _GEN_1119;
  wire [31:0] _GEN_1121 = 10'h79 == rs2[9:0] ? coeffs_121 : _GEN_1120;
  wire [31:0] _GEN_1122 = 10'h7a == rs2[9:0] ? coeffs_122 : _GEN_1121;
  wire [31:0] _GEN_1123 = 10'h7b == rs2[9:0] ? coeffs_123 : _GEN_1122;
  wire [31:0] _GEN_1124 = 10'h7c == rs2[9:0] ? coeffs_124 : _GEN_1123;
  wire [31:0] _GEN_1125 = 10'h7d == rs2[9:0] ? coeffs_125 : _GEN_1124;
  wire [31:0] _GEN_1126 = 10'h7e == rs2[9:0] ? coeffs_126 : _GEN_1125;
  wire [31:0] _GEN_1127 = 10'h7f == rs2[9:0] ? coeffs_127 : _GEN_1126;
  wire [31:0] _GEN_1128 = 10'h80 == rs2[9:0] ? coeffs_128 : _GEN_1127;
  wire [31:0] _GEN_1129 = 10'h81 == rs2[9:0] ? coeffs_129 : _GEN_1128;
  wire [31:0] _GEN_1130 = 10'h82 == rs2[9:0] ? coeffs_130 : _GEN_1129;
  wire [31:0] _GEN_1131 = 10'h83 == rs2[9:0] ? coeffs_131 : _GEN_1130;
  wire [31:0] _GEN_1132 = 10'h84 == rs2[9:0] ? coeffs_132 : _GEN_1131;
  wire [31:0] _GEN_1133 = 10'h85 == rs2[9:0] ? coeffs_133 : _GEN_1132;
  wire [31:0] _GEN_1134 = 10'h86 == rs2[9:0] ? coeffs_134 : _GEN_1133;
  wire [31:0] _GEN_1135 = 10'h87 == rs2[9:0] ? coeffs_135 : _GEN_1134;
  wire [31:0] _GEN_1136 = 10'h88 == rs2[9:0] ? coeffs_136 : _GEN_1135;
  wire [31:0] _GEN_1137 = 10'h89 == rs2[9:0] ? coeffs_137 : _GEN_1136;
  wire [31:0] _GEN_1138 = 10'h8a == rs2[9:0] ? coeffs_138 : _GEN_1137;
  wire [31:0] _GEN_1139 = 10'h8b == rs2[9:0] ? coeffs_139 : _GEN_1138;
  wire [31:0] _GEN_1140 = 10'h8c == rs2[9:0] ? coeffs_140 : _GEN_1139;
  wire [31:0] _GEN_1141 = 10'h8d == rs2[9:0] ? coeffs_141 : _GEN_1140;
  wire [31:0] _GEN_1142 = 10'h8e == rs2[9:0] ? coeffs_142 : _GEN_1141;
  wire [31:0] _GEN_1143 = 10'h8f == rs2[9:0] ? coeffs_143 : _GEN_1142;
  wire [31:0] _GEN_1144 = 10'h90 == rs2[9:0] ? coeffs_144 : _GEN_1143;
  wire [31:0] _GEN_1145 = 10'h91 == rs2[9:0] ? coeffs_145 : _GEN_1144;
  wire [31:0] _GEN_1146 = 10'h92 == rs2[9:0] ? coeffs_146 : _GEN_1145;
  wire [31:0] _GEN_1147 = 10'h93 == rs2[9:0] ? coeffs_147 : _GEN_1146;
  wire [31:0] _GEN_1148 = 10'h94 == rs2[9:0] ? coeffs_148 : _GEN_1147;
  wire [31:0] _GEN_1149 = 10'h95 == rs2[9:0] ? coeffs_149 : _GEN_1148;
  wire [31:0] _GEN_1150 = 10'h96 == rs2[9:0] ? coeffs_150 : _GEN_1149;
  wire [31:0] _GEN_1151 = 10'h97 == rs2[9:0] ? coeffs_151 : _GEN_1150;
  wire [31:0] _GEN_1152 = 10'h98 == rs2[9:0] ? coeffs_152 : _GEN_1151;
  wire [31:0] _GEN_1153 = 10'h99 == rs2[9:0] ? coeffs_153 : _GEN_1152;
  wire [31:0] _GEN_1154 = 10'h9a == rs2[9:0] ? coeffs_154 : _GEN_1153;
  wire [31:0] _GEN_1155 = 10'h9b == rs2[9:0] ? coeffs_155 : _GEN_1154;
  wire [31:0] _GEN_1156 = 10'h9c == rs2[9:0] ? coeffs_156 : _GEN_1155;
  wire [31:0] _GEN_1157 = 10'h9d == rs2[9:0] ? coeffs_157 : _GEN_1156;
  wire [31:0] _GEN_1158 = 10'h9e == rs2[9:0] ? coeffs_158 : _GEN_1157;
  wire [31:0] _GEN_1159 = 10'h9f == rs2[9:0] ? coeffs_159 : _GEN_1158;
  wire [31:0] _GEN_1160 = 10'ha0 == rs2[9:0] ? coeffs_160 : _GEN_1159;
  wire [31:0] _GEN_1161 = 10'ha1 == rs2[9:0] ? coeffs_161 : _GEN_1160;
  wire [31:0] _GEN_1162 = 10'ha2 == rs2[9:0] ? coeffs_162 : _GEN_1161;
  wire [31:0] _GEN_1163 = 10'ha3 == rs2[9:0] ? coeffs_163 : _GEN_1162;
  wire [31:0] _GEN_1164 = 10'ha4 == rs2[9:0] ? coeffs_164 : _GEN_1163;
  wire [31:0] _GEN_1165 = 10'ha5 == rs2[9:0] ? coeffs_165 : _GEN_1164;
  wire [31:0] _GEN_1166 = 10'ha6 == rs2[9:0] ? coeffs_166 : _GEN_1165;
  wire [31:0] _GEN_1167 = 10'ha7 == rs2[9:0] ? coeffs_167 : _GEN_1166;
  wire [31:0] _GEN_1168 = 10'ha8 == rs2[9:0] ? coeffs_168 : _GEN_1167;
  wire [31:0] _GEN_1169 = 10'ha9 == rs2[9:0] ? coeffs_169 : _GEN_1168;
  wire [31:0] _GEN_1170 = 10'haa == rs2[9:0] ? coeffs_170 : _GEN_1169;
  wire [31:0] _GEN_1171 = 10'hab == rs2[9:0] ? coeffs_171 : _GEN_1170;
  wire [31:0] _GEN_1172 = 10'hac == rs2[9:0] ? coeffs_172 : _GEN_1171;
  wire [31:0] _GEN_1173 = 10'had == rs2[9:0] ? coeffs_173 : _GEN_1172;
  wire [31:0] _GEN_1174 = 10'hae == rs2[9:0] ? coeffs_174 : _GEN_1173;
  wire [31:0] _GEN_1175 = 10'haf == rs2[9:0] ? coeffs_175 : _GEN_1174;
  wire [31:0] _GEN_1176 = 10'hb0 == rs2[9:0] ? coeffs_176 : _GEN_1175;
  wire [31:0] _GEN_1177 = 10'hb1 == rs2[9:0] ? coeffs_177 : _GEN_1176;
  wire [31:0] _GEN_1178 = 10'hb2 == rs2[9:0] ? coeffs_178 : _GEN_1177;
  wire [31:0] _GEN_1179 = 10'hb3 == rs2[9:0] ? coeffs_179 : _GEN_1178;
  wire [31:0] _GEN_1180 = 10'hb4 == rs2[9:0] ? coeffs_180 : _GEN_1179;
  wire [31:0] _GEN_1181 = 10'hb5 == rs2[9:0] ? coeffs_181 : _GEN_1180;
  wire [31:0] _GEN_1182 = 10'hb6 == rs2[9:0] ? coeffs_182 : _GEN_1181;
  wire [31:0] _GEN_1183 = 10'hb7 == rs2[9:0] ? coeffs_183 : _GEN_1182;
  wire [31:0] _GEN_1184 = 10'hb8 == rs2[9:0] ? coeffs_184 : _GEN_1183;
  wire [31:0] _GEN_1185 = 10'hb9 == rs2[9:0] ? coeffs_185 : _GEN_1184;
  wire [31:0] _GEN_1186 = 10'hba == rs2[9:0] ? coeffs_186 : _GEN_1185;
  wire [31:0] _GEN_1187 = 10'hbb == rs2[9:0] ? coeffs_187 : _GEN_1186;
  wire [31:0] _GEN_1188 = 10'hbc == rs2[9:0] ? coeffs_188 : _GEN_1187;
  wire [31:0] _GEN_1189 = 10'hbd == rs2[9:0] ? coeffs_189 : _GEN_1188;
  wire [31:0] _GEN_1190 = 10'hbe == rs2[9:0] ? coeffs_190 : _GEN_1189;
  wire [31:0] _GEN_1191 = 10'hbf == rs2[9:0] ? coeffs_191 : _GEN_1190;
  wire [31:0] _GEN_1192 = 10'hc0 == rs2[9:0] ? coeffs_192 : _GEN_1191;
  wire [31:0] _GEN_1193 = 10'hc1 == rs2[9:0] ? coeffs_193 : _GEN_1192;
  wire [31:0] _GEN_1194 = 10'hc2 == rs2[9:0] ? coeffs_194 : _GEN_1193;
  wire [31:0] _GEN_1195 = 10'hc3 == rs2[9:0] ? coeffs_195 : _GEN_1194;
  wire [31:0] _GEN_1196 = 10'hc4 == rs2[9:0] ? coeffs_196 : _GEN_1195;
  wire [31:0] _GEN_1197 = 10'hc5 == rs2[9:0] ? coeffs_197 : _GEN_1196;
  wire [31:0] _GEN_1198 = 10'hc6 == rs2[9:0] ? coeffs_198 : _GEN_1197;
  wire [31:0] _GEN_1199 = 10'hc7 == rs2[9:0] ? coeffs_199 : _GEN_1198;
  wire [31:0] _GEN_1200 = 10'hc8 == rs2[9:0] ? coeffs_200 : _GEN_1199;
  wire [31:0] _GEN_1201 = 10'hc9 == rs2[9:0] ? coeffs_201 : _GEN_1200;
  wire [31:0] _GEN_1202 = 10'hca == rs2[9:0] ? coeffs_202 : _GEN_1201;
  wire [31:0] _GEN_1203 = 10'hcb == rs2[9:0] ? coeffs_203 : _GEN_1202;
  wire [31:0] _GEN_1204 = 10'hcc == rs2[9:0] ? coeffs_204 : _GEN_1203;
  wire [31:0] _GEN_1205 = 10'hcd == rs2[9:0] ? coeffs_205 : _GEN_1204;
  wire [31:0] _GEN_1206 = 10'hce == rs2[9:0] ? coeffs_206 : _GEN_1205;
  wire [31:0] _GEN_1207 = 10'hcf == rs2[9:0] ? coeffs_207 : _GEN_1206;
  wire [31:0] _GEN_1208 = 10'hd0 == rs2[9:0] ? coeffs_208 : _GEN_1207;
  wire [31:0] _GEN_1209 = 10'hd1 == rs2[9:0] ? coeffs_209 : _GEN_1208;
  wire [31:0] _GEN_1210 = 10'hd2 == rs2[9:0] ? coeffs_210 : _GEN_1209;
  wire [31:0] _GEN_1211 = 10'hd3 == rs2[9:0] ? coeffs_211 : _GEN_1210;
  wire [31:0] _GEN_1212 = 10'hd4 == rs2[9:0] ? coeffs_212 : _GEN_1211;
  wire [31:0] _GEN_1213 = 10'hd5 == rs2[9:0] ? coeffs_213 : _GEN_1212;
  wire [31:0] _GEN_1214 = 10'hd6 == rs2[9:0] ? coeffs_214 : _GEN_1213;
  wire [31:0] _GEN_1215 = 10'hd7 == rs2[9:0] ? coeffs_215 : _GEN_1214;
  wire [31:0] _GEN_1216 = 10'hd8 == rs2[9:0] ? coeffs_216 : _GEN_1215;
  wire [31:0] _GEN_1217 = 10'hd9 == rs2[9:0] ? coeffs_217 : _GEN_1216;
  wire [31:0] _GEN_1218 = 10'hda == rs2[9:0] ? coeffs_218 : _GEN_1217;
  wire [31:0] _GEN_1219 = 10'hdb == rs2[9:0] ? coeffs_219 : _GEN_1218;
  wire [31:0] _GEN_1220 = 10'hdc == rs2[9:0] ? coeffs_220 : _GEN_1219;
  wire [31:0] _GEN_1221 = 10'hdd == rs2[9:0] ? coeffs_221 : _GEN_1220;
  wire [31:0] _GEN_1222 = 10'hde == rs2[9:0] ? coeffs_222 : _GEN_1221;
  wire [31:0] _GEN_1223 = 10'hdf == rs2[9:0] ? coeffs_223 : _GEN_1222;
  wire [31:0] _GEN_1224 = 10'he0 == rs2[9:0] ? coeffs_224 : _GEN_1223;
  wire [31:0] _GEN_1225 = 10'he1 == rs2[9:0] ? coeffs_225 : _GEN_1224;
  wire [31:0] _GEN_1226 = 10'he2 == rs2[9:0] ? coeffs_226 : _GEN_1225;
  wire [31:0] _GEN_1227 = 10'he3 == rs2[9:0] ? coeffs_227 : _GEN_1226;
  wire [31:0] _GEN_1228 = 10'he4 == rs2[9:0] ? coeffs_228 : _GEN_1227;
  wire [31:0] _GEN_1229 = 10'he5 == rs2[9:0] ? coeffs_229 : _GEN_1228;
  wire [31:0] _GEN_1230 = 10'he6 == rs2[9:0] ? coeffs_230 : _GEN_1229;
  wire [31:0] _GEN_1231 = 10'he7 == rs2[9:0] ? coeffs_231 : _GEN_1230;
  wire [31:0] _GEN_1232 = 10'he8 == rs2[9:0] ? coeffs_232 : _GEN_1231;
  wire [31:0] _GEN_1233 = 10'he9 == rs2[9:0] ? coeffs_233 : _GEN_1232;
  wire [31:0] _GEN_1234 = 10'hea == rs2[9:0] ? coeffs_234 : _GEN_1233;
  wire [31:0] _GEN_1235 = 10'heb == rs2[9:0] ? coeffs_235 : _GEN_1234;
  wire [31:0] _GEN_1236 = 10'hec == rs2[9:0] ? coeffs_236 : _GEN_1235;
  wire [31:0] _GEN_1237 = 10'hed == rs2[9:0] ? coeffs_237 : _GEN_1236;
  wire [31:0] _GEN_1238 = 10'hee == rs2[9:0] ? coeffs_238 : _GEN_1237;
  wire [31:0] _GEN_1239 = 10'hef == rs2[9:0] ? coeffs_239 : _GEN_1238;
  wire [31:0] _GEN_1240 = 10'hf0 == rs2[9:0] ? coeffs_240 : _GEN_1239;
  wire [31:0] _GEN_1241 = 10'hf1 == rs2[9:0] ? coeffs_241 : _GEN_1240;
  wire [31:0] _GEN_1242 = 10'hf2 == rs2[9:0] ? coeffs_242 : _GEN_1241;
  wire [31:0] _GEN_1243 = 10'hf3 == rs2[9:0] ? coeffs_243 : _GEN_1242;
  wire [31:0] _GEN_1244 = 10'hf4 == rs2[9:0] ? coeffs_244 : _GEN_1243;
  wire [31:0] _GEN_1245 = 10'hf5 == rs2[9:0] ? coeffs_245 : _GEN_1244;
  wire [31:0] _GEN_1246 = 10'hf6 == rs2[9:0] ? coeffs_246 : _GEN_1245;
  wire [31:0] _GEN_1247 = 10'hf7 == rs2[9:0] ? coeffs_247 : _GEN_1246;
  wire [31:0] _GEN_1248 = 10'hf8 == rs2[9:0] ? coeffs_248 : _GEN_1247;
  wire [31:0] _GEN_1249 = 10'hf9 == rs2[9:0] ? coeffs_249 : _GEN_1248;
  wire [31:0] _GEN_1250 = 10'hfa == rs2[9:0] ? coeffs_250 : _GEN_1249;
  wire [31:0] _GEN_1251 = 10'hfb == rs2[9:0] ? coeffs_251 : _GEN_1250;
  wire [31:0] _GEN_1252 = 10'hfc == rs2[9:0] ? coeffs_252 : _GEN_1251;
  wire [31:0] _GEN_1253 = 10'hfd == rs2[9:0] ? coeffs_253 : _GEN_1252;
  wire [31:0] _GEN_1254 = 10'hfe == rs2[9:0] ? coeffs_254 : _GEN_1253;
  wire [31:0] _GEN_1255 = 10'hff == rs2[9:0] ? coeffs_255 : _GEN_1254;
  wire [31:0] _GEN_1256 = 10'h100 == rs2[9:0] ? coeffs_256 : _GEN_1255;
  wire [31:0] _GEN_1257 = 10'h101 == rs2[9:0] ? coeffs_257 : _GEN_1256;
  wire [31:0] _GEN_1258 = 10'h102 == rs2[9:0] ? coeffs_258 : _GEN_1257;
  wire [31:0] _GEN_1259 = 10'h103 == rs2[9:0] ? coeffs_259 : _GEN_1258;
  wire [31:0] _GEN_1260 = 10'h104 == rs2[9:0] ? coeffs_260 : _GEN_1259;
  wire [31:0] _GEN_1261 = 10'h105 == rs2[9:0] ? coeffs_261 : _GEN_1260;
  wire [31:0] _GEN_1262 = 10'h106 == rs2[9:0] ? coeffs_262 : _GEN_1261;
  wire [31:0] _GEN_1263 = 10'h107 == rs2[9:0] ? coeffs_263 : _GEN_1262;
  wire [31:0] _GEN_1264 = 10'h108 == rs2[9:0] ? coeffs_264 : _GEN_1263;
  wire [31:0] _GEN_1265 = 10'h109 == rs2[9:0] ? coeffs_265 : _GEN_1264;
  wire [31:0] _GEN_1266 = 10'h10a == rs2[9:0] ? coeffs_266 : _GEN_1265;
  wire [31:0] _GEN_1267 = 10'h10b == rs2[9:0] ? coeffs_267 : _GEN_1266;
  wire [31:0] _GEN_1268 = 10'h10c == rs2[9:0] ? coeffs_268 : _GEN_1267;
  wire [31:0] _GEN_1269 = 10'h10d == rs2[9:0] ? coeffs_269 : _GEN_1268;
  wire [31:0] _GEN_1270 = 10'h10e == rs2[9:0] ? coeffs_270 : _GEN_1269;
  wire [31:0] _GEN_1271 = 10'h10f == rs2[9:0] ? coeffs_271 : _GEN_1270;
  wire [31:0] _GEN_1272 = 10'h110 == rs2[9:0] ? coeffs_272 : _GEN_1271;
  wire [31:0] _GEN_1273 = 10'h111 == rs2[9:0] ? coeffs_273 : _GEN_1272;
  wire [31:0] _GEN_1274 = 10'h112 == rs2[9:0] ? coeffs_274 : _GEN_1273;
  wire [31:0] _GEN_1275 = 10'h113 == rs2[9:0] ? coeffs_275 : _GEN_1274;
  wire [31:0] _GEN_1276 = 10'h114 == rs2[9:0] ? coeffs_276 : _GEN_1275;
  wire [31:0] _GEN_1277 = 10'h115 == rs2[9:0] ? coeffs_277 : _GEN_1276;
  wire [31:0] _GEN_1278 = 10'h116 == rs2[9:0] ? coeffs_278 : _GEN_1277;
  wire [31:0] _GEN_1279 = 10'h117 == rs2[9:0] ? coeffs_279 : _GEN_1278;
  wire [31:0] _GEN_1280 = 10'h118 == rs2[9:0] ? coeffs_280 : _GEN_1279;
  wire [31:0] _GEN_1281 = 10'h119 == rs2[9:0] ? coeffs_281 : _GEN_1280;
  wire [31:0] _GEN_1282 = 10'h11a == rs2[9:0] ? coeffs_282 : _GEN_1281;
  wire [31:0] _GEN_1283 = 10'h11b == rs2[9:0] ? coeffs_283 : _GEN_1282;
  wire [31:0] _GEN_1284 = 10'h11c == rs2[9:0] ? coeffs_284 : _GEN_1283;
  wire [31:0] _GEN_1285 = 10'h11d == rs2[9:0] ? coeffs_285 : _GEN_1284;
  wire [31:0] _GEN_1286 = 10'h11e == rs2[9:0] ? coeffs_286 : _GEN_1285;
  wire [31:0] _GEN_1287 = 10'h11f == rs2[9:0] ? coeffs_287 : _GEN_1286;
  wire [31:0] _GEN_1288 = 10'h120 == rs2[9:0] ? coeffs_288 : _GEN_1287;
  wire [31:0] _GEN_1289 = 10'h121 == rs2[9:0] ? coeffs_289 : _GEN_1288;
  wire [31:0] _GEN_1290 = 10'h122 == rs2[9:0] ? coeffs_290 : _GEN_1289;
  wire [31:0] _GEN_1291 = 10'h123 == rs2[9:0] ? coeffs_291 : _GEN_1290;
  wire [31:0] _GEN_1292 = 10'h124 == rs2[9:0] ? coeffs_292 : _GEN_1291;
  wire [31:0] _GEN_1293 = 10'h125 == rs2[9:0] ? coeffs_293 : _GEN_1292;
  wire [31:0] _GEN_1294 = 10'h126 == rs2[9:0] ? coeffs_294 : _GEN_1293;
  wire [31:0] _GEN_1295 = 10'h127 == rs2[9:0] ? coeffs_295 : _GEN_1294;
  wire [31:0] _GEN_1296 = 10'h128 == rs2[9:0] ? coeffs_296 : _GEN_1295;
  wire [31:0] _GEN_1297 = 10'h129 == rs2[9:0] ? coeffs_297 : _GEN_1296;
  wire [31:0] _GEN_1298 = 10'h12a == rs2[9:0] ? coeffs_298 : _GEN_1297;
  wire [31:0] _GEN_1299 = 10'h12b == rs2[9:0] ? coeffs_299 : _GEN_1298;
  wire [31:0] _GEN_1300 = 10'h12c == rs2[9:0] ? coeffs_300 : _GEN_1299;
  wire [31:0] _GEN_1301 = 10'h12d == rs2[9:0] ? coeffs_301 : _GEN_1300;
  wire [31:0] _GEN_1302 = 10'h12e == rs2[9:0] ? coeffs_302 : _GEN_1301;
  wire [31:0] _GEN_1303 = 10'h12f == rs2[9:0] ? coeffs_303 : _GEN_1302;
  wire [31:0] _GEN_1304 = 10'h130 == rs2[9:0] ? coeffs_304 : _GEN_1303;
  wire [31:0] _GEN_1305 = 10'h131 == rs2[9:0] ? coeffs_305 : _GEN_1304;
  wire [31:0] _GEN_1306 = 10'h132 == rs2[9:0] ? coeffs_306 : _GEN_1305;
  wire [31:0] _GEN_1307 = 10'h133 == rs2[9:0] ? coeffs_307 : _GEN_1306;
  wire [31:0] _GEN_1308 = 10'h134 == rs2[9:0] ? coeffs_308 : _GEN_1307;
  wire [31:0] _GEN_1309 = 10'h135 == rs2[9:0] ? coeffs_309 : _GEN_1308;
  wire [31:0] _GEN_1310 = 10'h136 == rs2[9:0] ? coeffs_310 : _GEN_1309;
  wire [31:0] _GEN_1311 = 10'h137 == rs2[9:0] ? coeffs_311 : _GEN_1310;
  wire [31:0] _GEN_1312 = 10'h138 == rs2[9:0] ? coeffs_312 : _GEN_1311;
  wire [31:0] _GEN_1313 = 10'h139 == rs2[9:0] ? coeffs_313 : _GEN_1312;
  wire [31:0] _GEN_1314 = 10'h13a == rs2[9:0] ? coeffs_314 : _GEN_1313;
  wire [31:0] _GEN_1315 = 10'h13b == rs2[9:0] ? coeffs_315 : _GEN_1314;
  wire [31:0] _GEN_1316 = 10'h13c == rs2[9:0] ? coeffs_316 : _GEN_1315;
  wire [31:0] _GEN_1317 = 10'h13d == rs2[9:0] ? coeffs_317 : _GEN_1316;
  wire [31:0] _GEN_1318 = 10'h13e == rs2[9:0] ? coeffs_318 : _GEN_1317;
  wire [31:0] _GEN_1319 = 10'h13f == rs2[9:0] ? coeffs_319 : _GEN_1318;
  wire [31:0] _GEN_1320 = 10'h140 == rs2[9:0] ? coeffs_320 : _GEN_1319;
  wire [31:0] _GEN_1321 = 10'h141 == rs2[9:0] ? coeffs_321 : _GEN_1320;
  wire [31:0] _GEN_1322 = 10'h142 == rs2[9:0] ? coeffs_322 : _GEN_1321;
  wire [31:0] _GEN_1323 = 10'h143 == rs2[9:0] ? coeffs_323 : _GEN_1322;
  wire [31:0] _GEN_1324 = 10'h144 == rs2[9:0] ? coeffs_324 : _GEN_1323;
  wire [31:0] _GEN_1325 = 10'h145 == rs2[9:0] ? coeffs_325 : _GEN_1324;
  wire [31:0] _GEN_1326 = 10'h146 == rs2[9:0] ? coeffs_326 : _GEN_1325;
  wire [31:0] _GEN_1327 = 10'h147 == rs2[9:0] ? coeffs_327 : _GEN_1326;
  wire [31:0] _GEN_1328 = 10'h148 == rs2[9:0] ? coeffs_328 : _GEN_1327;
  wire [31:0] _GEN_1329 = 10'h149 == rs2[9:0] ? coeffs_329 : _GEN_1328;
  wire [31:0] _GEN_1330 = 10'h14a == rs2[9:0] ? coeffs_330 : _GEN_1329;
  wire [31:0] _GEN_1331 = 10'h14b == rs2[9:0] ? coeffs_331 : _GEN_1330;
  wire [31:0] _GEN_1332 = 10'h14c == rs2[9:0] ? coeffs_332 : _GEN_1331;
  wire [31:0] _GEN_1333 = 10'h14d == rs2[9:0] ? coeffs_333 : _GEN_1332;
  wire [31:0] _GEN_1334 = 10'h14e == rs2[9:0] ? coeffs_334 : _GEN_1333;
  wire [31:0] _GEN_1335 = 10'h14f == rs2[9:0] ? coeffs_335 : _GEN_1334;
  wire [31:0] _GEN_1336 = 10'h150 == rs2[9:0] ? coeffs_336 : _GEN_1335;
  wire [31:0] _GEN_1337 = 10'h151 == rs2[9:0] ? coeffs_337 : _GEN_1336;
  wire [31:0] _GEN_1338 = 10'h152 == rs2[9:0] ? coeffs_338 : _GEN_1337;
  wire [31:0] _GEN_1339 = 10'h153 == rs2[9:0] ? coeffs_339 : _GEN_1338;
  wire [31:0] _GEN_1340 = 10'h154 == rs2[9:0] ? coeffs_340 : _GEN_1339;
  wire [31:0] _GEN_1341 = 10'h155 == rs2[9:0] ? coeffs_341 : _GEN_1340;
  wire [31:0] _GEN_1342 = 10'h156 == rs2[9:0] ? coeffs_342 : _GEN_1341;
  wire [31:0] _GEN_1343 = 10'h157 == rs2[9:0] ? coeffs_343 : _GEN_1342;
  wire [31:0] _GEN_1344 = 10'h158 == rs2[9:0] ? coeffs_344 : _GEN_1343;
  wire [31:0] _GEN_1345 = 10'h159 == rs2[9:0] ? coeffs_345 : _GEN_1344;
  wire [31:0] _GEN_1346 = 10'h15a == rs2[9:0] ? coeffs_346 : _GEN_1345;
  wire [31:0] _GEN_1347 = 10'h15b == rs2[9:0] ? coeffs_347 : _GEN_1346;
  wire [31:0] _GEN_1348 = 10'h15c == rs2[9:0] ? coeffs_348 : _GEN_1347;
  wire [31:0] _GEN_1349 = 10'h15d == rs2[9:0] ? coeffs_349 : _GEN_1348;
  wire [31:0] _GEN_1350 = 10'h15e == rs2[9:0] ? coeffs_350 : _GEN_1349;
  wire [31:0] _GEN_1351 = 10'h15f == rs2[9:0] ? coeffs_351 : _GEN_1350;
  wire [31:0] _GEN_1352 = 10'h160 == rs2[9:0] ? coeffs_352 : _GEN_1351;
  wire [31:0] _GEN_1353 = 10'h161 == rs2[9:0] ? coeffs_353 : _GEN_1352;
  wire [31:0] _GEN_1354 = 10'h162 == rs2[9:0] ? coeffs_354 : _GEN_1353;
  wire [31:0] _GEN_1355 = 10'h163 == rs2[9:0] ? coeffs_355 : _GEN_1354;
  wire [31:0] _GEN_1356 = 10'h164 == rs2[9:0] ? coeffs_356 : _GEN_1355;
  wire [31:0] _GEN_1357 = 10'h165 == rs2[9:0] ? coeffs_357 : _GEN_1356;
  wire [31:0] _GEN_1358 = 10'h166 == rs2[9:0] ? coeffs_358 : _GEN_1357;
  wire [31:0] _GEN_1359 = 10'h167 == rs2[9:0] ? coeffs_359 : _GEN_1358;
  wire [31:0] _GEN_1360 = 10'h168 == rs2[9:0] ? coeffs_360 : _GEN_1359;
  wire [31:0] _GEN_1361 = 10'h169 == rs2[9:0] ? coeffs_361 : _GEN_1360;
  wire [31:0] _GEN_1362 = 10'h16a == rs2[9:0] ? coeffs_362 : _GEN_1361;
  wire [31:0] _GEN_1363 = 10'h16b == rs2[9:0] ? coeffs_363 : _GEN_1362;
  wire [31:0] _GEN_1364 = 10'h16c == rs2[9:0] ? coeffs_364 : _GEN_1363;
  wire [31:0] _GEN_1365 = 10'h16d == rs2[9:0] ? coeffs_365 : _GEN_1364;
  wire [31:0] _GEN_1366 = 10'h16e == rs2[9:0] ? coeffs_366 : _GEN_1365;
  wire [31:0] _GEN_1367 = 10'h16f == rs2[9:0] ? coeffs_367 : _GEN_1366;
  wire [31:0] _GEN_1368 = 10'h170 == rs2[9:0] ? coeffs_368 : _GEN_1367;
  wire [31:0] _GEN_1369 = 10'h171 == rs2[9:0] ? coeffs_369 : _GEN_1368;
  wire [31:0] _GEN_1370 = 10'h172 == rs2[9:0] ? coeffs_370 : _GEN_1369;
  wire [31:0] _GEN_1371 = 10'h173 == rs2[9:0] ? coeffs_371 : _GEN_1370;
  wire [31:0] _GEN_1372 = 10'h174 == rs2[9:0] ? coeffs_372 : _GEN_1371;
  wire [31:0] _GEN_1373 = 10'h175 == rs2[9:0] ? coeffs_373 : _GEN_1372;
  wire [31:0] _GEN_1374 = 10'h176 == rs2[9:0] ? coeffs_374 : _GEN_1373;
  wire [31:0] _GEN_1375 = 10'h177 == rs2[9:0] ? coeffs_375 : _GEN_1374;
  wire [31:0] _GEN_1376 = 10'h178 == rs2[9:0] ? coeffs_376 : _GEN_1375;
  wire [31:0] _GEN_1377 = 10'h179 == rs2[9:0] ? coeffs_377 : _GEN_1376;
  wire [31:0] _GEN_1378 = 10'h17a == rs2[9:0] ? coeffs_378 : _GEN_1377;
  wire [31:0] _GEN_1379 = 10'h17b == rs2[9:0] ? coeffs_379 : _GEN_1378;
  wire [31:0] _GEN_1380 = 10'h17c == rs2[9:0] ? coeffs_380 : _GEN_1379;
  wire [31:0] _GEN_1381 = 10'h17d == rs2[9:0] ? coeffs_381 : _GEN_1380;
  wire [31:0] _GEN_1382 = 10'h17e == rs2[9:0] ? coeffs_382 : _GEN_1381;
  wire [31:0] _GEN_1383 = 10'h17f == rs2[9:0] ? coeffs_383 : _GEN_1382;
  wire [31:0] _GEN_1384 = 10'h180 == rs2[9:0] ? coeffs_384 : _GEN_1383;
  wire [31:0] _GEN_1385 = 10'h181 == rs2[9:0] ? coeffs_385 : _GEN_1384;
  wire [31:0] _GEN_1386 = 10'h182 == rs2[9:0] ? coeffs_386 : _GEN_1385;
  wire [31:0] _GEN_1387 = 10'h183 == rs2[9:0] ? coeffs_387 : _GEN_1386;
  wire [31:0] _GEN_1388 = 10'h184 == rs2[9:0] ? coeffs_388 : _GEN_1387;
  wire [31:0] _GEN_1389 = 10'h185 == rs2[9:0] ? coeffs_389 : _GEN_1388;
  wire [31:0] _GEN_1390 = 10'h186 == rs2[9:0] ? coeffs_390 : _GEN_1389;
  wire [31:0] _GEN_1391 = 10'h187 == rs2[9:0] ? coeffs_391 : _GEN_1390;
  wire [31:0] _GEN_1392 = 10'h188 == rs2[9:0] ? coeffs_392 : _GEN_1391;
  wire [31:0] _GEN_1393 = 10'h189 == rs2[9:0] ? coeffs_393 : _GEN_1392;
  wire [31:0] _GEN_1394 = 10'h18a == rs2[9:0] ? coeffs_394 : _GEN_1393;
  wire [31:0] _GEN_1395 = 10'h18b == rs2[9:0] ? coeffs_395 : _GEN_1394;
  wire [31:0] _GEN_1396 = 10'h18c == rs2[9:0] ? coeffs_396 : _GEN_1395;
  wire [31:0] _GEN_1397 = 10'h18d == rs2[9:0] ? coeffs_397 : _GEN_1396;
  wire [31:0] _GEN_1398 = 10'h18e == rs2[9:0] ? coeffs_398 : _GEN_1397;
  wire [31:0] _GEN_1399 = 10'h18f == rs2[9:0] ? coeffs_399 : _GEN_1398;
  wire [31:0] _GEN_1400 = 10'h190 == rs2[9:0] ? coeffs_400 : _GEN_1399;
  wire [31:0] _GEN_1401 = 10'h191 == rs2[9:0] ? coeffs_401 : _GEN_1400;
  wire [31:0] _GEN_1402 = 10'h192 == rs2[9:0] ? coeffs_402 : _GEN_1401;
  wire [31:0] _GEN_1403 = 10'h193 == rs2[9:0] ? coeffs_403 : _GEN_1402;
  wire [31:0] _GEN_1404 = 10'h194 == rs2[9:0] ? coeffs_404 : _GEN_1403;
  wire [31:0] _GEN_1405 = 10'h195 == rs2[9:0] ? coeffs_405 : _GEN_1404;
  wire [31:0] _GEN_1406 = 10'h196 == rs2[9:0] ? coeffs_406 : _GEN_1405;
  wire [31:0] _GEN_1407 = 10'h197 == rs2[9:0] ? coeffs_407 : _GEN_1406;
  wire [31:0] _GEN_1408 = 10'h198 == rs2[9:0] ? coeffs_408 : _GEN_1407;
  wire [31:0] _GEN_1409 = 10'h199 == rs2[9:0] ? coeffs_409 : _GEN_1408;
  wire [31:0] _GEN_1410 = 10'h19a == rs2[9:0] ? coeffs_410 : _GEN_1409;
  wire [31:0] _GEN_1411 = 10'h19b == rs2[9:0] ? coeffs_411 : _GEN_1410;
  wire [31:0] _GEN_1412 = 10'h19c == rs2[9:0] ? coeffs_412 : _GEN_1411;
  wire [31:0] _GEN_1413 = 10'h19d == rs2[9:0] ? coeffs_413 : _GEN_1412;
  wire [31:0] _GEN_1414 = 10'h19e == rs2[9:0] ? coeffs_414 : _GEN_1413;
  wire [31:0] _GEN_1415 = 10'h19f == rs2[9:0] ? coeffs_415 : _GEN_1414;
  wire [31:0] _GEN_1416 = 10'h1a0 == rs2[9:0] ? coeffs_416 : _GEN_1415;
  wire [31:0] _GEN_1417 = 10'h1a1 == rs2[9:0] ? coeffs_417 : _GEN_1416;
  wire [31:0] _GEN_1418 = 10'h1a2 == rs2[9:0] ? coeffs_418 : _GEN_1417;
  wire [31:0] _GEN_1419 = 10'h1a3 == rs2[9:0] ? coeffs_419 : _GEN_1418;
  wire [31:0] _GEN_1420 = 10'h1a4 == rs2[9:0] ? coeffs_420 : _GEN_1419;
  wire [31:0] _GEN_1421 = 10'h1a5 == rs2[9:0] ? coeffs_421 : _GEN_1420;
  wire [31:0] _GEN_1422 = 10'h1a6 == rs2[9:0] ? coeffs_422 : _GEN_1421;
  wire [31:0] _GEN_1423 = 10'h1a7 == rs2[9:0] ? coeffs_423 : _GEN_1422;
  wire [31:0] _GEN_1424 = 10'h1a8 == rs2[9:0] ? coeffs_424 : _GEN_1423;
  wire [31:0] _GEN_1425 = 10'h1a9 == rs2[9:0] ? coeffs_425 : _GEN_1424;
  wire [31:0] _GEN_1426 = 10'h1aa == rs2[9:0] ? coeffs_426 : _GEN_1425;
  wire [31:0] _GEN_1427 = 10'h1ab == rs2[9:0] ? coeffs_427 : _GEN_1426;
  wire [31:0] _GEN_1428 = 10'h1ac == rs2[9:0] ? coeffs_428 : _GEN_1427;
  wire [31:0] _GEN_1429 = 10'h1ad == rs2[9:0] ? coeffs_429 : _GEN_1428;
  wire [31:0] _GEN_1430 = 10'h1ae == rs2[9:0] ? coeffs_430 : _GEN_1429;
  wire [31:0] _GEN_1431 = 10'h1af == rs2[9:0] ? coeffs_431 : _GEN_1430;
  wire [31:0] _GEN_1432 = 10'h1b0 == rs2[9:0] ? coeffs_432 : _GEN_1431;
  wire [31:0] _GEN_1433 = 10'h1b1 == rs2[9:0] ? coeffs_433 : _GEN_1432;
  wire [31:0] _GEN_1434 = 10'h1b2 == rs2[9:0] ? coeffs_434 : _GEN_1433;
  wire [31:0] _GEN_1435 = 10'h1b3 == rs2[9:0] ? coeffs_435 : _GEN_1434;
  wire [31:0] _GEN_1436 = 10'h1b4 == rs2[9:0] ? coeffs_436 : _GEN_1435;
  wire [31:0] _GEN_1437 = 10'h1b5 == rs2[9:0] ? coeffs_437 : _GEN_1436;
  wire [31:0] _GEN_1438 = 10'h1b6 == rs2[9:0] ? coeffs_438 : _GEN_1437;
  wire [31:0] _GEN_1439 = 10'h1b7 == rs2[9:0] ? coeffs_439 : _GEN_1438;
  wire [31:0] _GEN_1440 = 10'h1b8 == rs2[9:0] ? coeffs_440 : _GEN_1439;
  wire [31:0] _GEN_1441 = 10'h1b9 == rs2[9:0] ? coeffs_441 : _GEN_1440;
  wire [31:0] _GEN_1442 = 10'h1ba == rs2[9:0] ? coeffs_442 : _GEN_1441;
  wire [31:0] _GEN_1443 = 10'h1bb == rs2[9:0] ? coeffs_443 : _GEN_1442;
  wire [31:0] _GEN_1444 = 10'h1bc == rs2[9:0] ? coeffs_444 : _GEN_1443;
  wire [31:0] _GEN_1445 = 10'h1bd == rs2[9:0] ? coeffs_445 : _GEN_1444;
  wire [31:0] _GEN_1446 = 10'h1be == rs2[9:0] ? coeffs_446 : _GEN_1445;
  wire [31:0] _GEN_1447 = 10'h1bf == rs2[9:0] ? coeffs_447 : _GEN_1446;
  wire [31:0] _GEN_1448 = 10'h1c0 == rs2[9:0] ? coeffs_448 : _GEN_1447;
  wire [31:0] _GEN_1449 = 10'h1c1 == rs2[9:0] ? coeffs_449 : _GEN_1448;
  wire [31:0] _GEN_1450 = 10'h1c2 == rs2[9:0] ? coeffs_450 : _GEN_1449;
  wire [31:0] _GEN_1451 = 10'h1c3 == rs2[9:0] ? coeffs_451 : _GEN_1450;
  wire [31:0] _GEN_1452 = 10'h1c4 == rs2[9:0] ? coeffs_452 : _GEN_1451;
  wire [31:0] _GEN_1453 = 10'h1c5 == rs2[9:0] ? coeffs_453 : _GEN_1452;
  wire [31:0] _GEN_1454 = 10'h1c6 == rs2[9:0] ? coeffs_454 : _GEN_1453;
  wire [31:0] _GEN_1455 = 10'h1c7 == rs2[9:0] ? coeffs_455 : _GEN_1454;
  wire [31:0] _GEN_1456 = 10'h1c8 == rs2[9:0] ? coeffs_456 : _GEN_1455;
  wire [31:0] _GEN_1457 = 10'h1c9 == rs2[9:0] ? coeffs_457 : _GEN_1456;
  wire [31:0] _GEN_1458 = 10'h1ca == rs2[9:0] ? coeffs_458 : _GEN_1457;
  wire [31:0] _GEN_1459 = 10'h1cb == rs2[9:0] ? coeffs_459 : _GEN_1458;
  wire [31:0] _GEN_1460 = 10'h1cc == rs2[9:0] ? coeffs_460 : _GEN_1459;
  wire [31:0] _GEN_1461 = 10'h1cd == rs2[9:0] ? coeffs_461 : _GEN_1460;
  wire [31:0] _GEN_1462 = 10'h1ce == rs2[9:0] ? coeffs_462 : _GEN_1461;
  wire [31:0] _GEN_1463 = 10'h1cf == rs2[9:0] ? coeffs_463 : _GEN_1462;
  wire [31:0] _GEN_1464 = 10'h1d0 == rs2[9:0] ? coeffs_464 : _GEN_1463;
  wire [31:0] _GEN_1465 = 10'h1d1 == rs2[9:0] ? coeffs_465 : _GEN_1464;
  wire [31:0] _GEN_1466 = 10'h1d2 == rs2[9:0] ? coeffs_466 : _GEN_1465;
  wire [31:0] _GEN_1467 = 10'h1d3 == rs2[9:0] ? coeffs_467 : _GEN_1466;
  wire [31:0] _GEN_1468 = 10'h1d4 == rs2[9:0] ? coeffs_468 : _GEN_1467;
  wire [31:0] _GEN_1469 = 10'h1d5 == rs2[9:0] ? coeffs_469 : _GEN_1468;
  wire [31:0] _GEN_1470 = 10'h1d6 == rs2[9:0] ? coeffs_470 : _GEN_1469;
  wire [31:0] _GEN_1471 = 10'h1d7 == rs2[9:0] ? coeffs_471 : _GEN_1470;
  wire [31:0] _GEN_1472 = 10'h1d8 == rs2[9:0] ? coeffs_472 : _GEN_1471;
  wire [31:0] _GEN_1473 = 10'h1d9 == rs2[9:0] ? coeffs_473 : _GEN_1472;
  wire [31:0] _GEN_1474 = 10'h1da == rs2[9:0] ? coeffs_474 : _GEN_1473;
  wire [31:0] _GEN_1475 = 10'h1db == rs2[9:0] ? coeffs_475 : _GEN_1474;
  wire [31:0] _GEN_1476 = 10'h1dc == rs2[9:0] ? coeffs_476 : _GEN_1475;
  wire [31:0] _GEN_1477 = 10'h1dd == rs2[9:0] ? coeffs_477 : _GEN_1476;
  wire [31:0] _GEN_1478 = 10'h1de == rs2[9:0] ? coeffs_478 : _GEN_1477;
  wire [31:0] _GEN_1479 = 10'h1df == rs2[9:0] ? coeffs_479 : _GEN_1478;
  wire [31:0] _GEN_1480 = 10'h1e0 == rs2[9:0] ? coeffs_480 : _GEN_1479;
  wire [31:0] _GEN_1481 = 10'h1e1 == rs2[9:0] ? coeffs_481 : _GEN_1480;
  wire [31:0] _GEN_1482 = 10'h1e2 == rs2[9:0] ? coeffs_482 : _GEN_1481;
  wire [31:0] _GEN_1483 = 10'h1e3 == rs2[9:0] ? coeffs_483 : _GEN_1482;
  wire [31:0] _GEN_1484 = 10'h1e4 == rs2[9:0] ? coeffs_484 : _GEN_1483;
  wire [31:0] _GEN_1485 = 10'h1e5 == rs2[9:0] ? coeffs_485 : _GEN_1484;
  wire [31:0] _GEN_1486 = 10'h1e6 == rs2[9:0] ? coeffs_486 : _GEN_1485;
  wire [31:0] _GEN_1487 = 10'h1e7 == rs2[9:0] ? coeffs_487 : _GEN_1486;
  wire [31:0] _GEN_1488 = 10'h1e8 == rs2[9:0] ? coeffs_488 : _GEN_1487;
  wire [31:0] _GEN_1489 = 10'h1e9 == rs2[9:0] ? coeffs_489 : _GEN_1488;
  wire [31:0] _GEN_1490 = 10'h1ea == rs2[9:0] ? coeffs_490 : _GEN_1489;
  wire [31:0] _GEN_1491 = 10'h1eb == rs2[9:0] ? coeffs_491 : _GEN_1490;
  wire [31:0] _GEN_1492 = 10'h1ec == rs2[9:0] ? coeffs_492 : _GEN_1491;
  wire [31:0] _GEN_1493 = 10'h1ed == rs2[9:0] ? coeffs_493 : _GEN_1492;
  wire [31:0] _GEN_1494 = 10'h1ee == rs2[9:0] ? coeffs_494 : _GEN_1493;
  wire [31:0] _GEN_1495 = 10'h1ef == rs2[9:0] ? coeffs_495 : _GEN_1494;
  wire [31:0] _GEN_1496 = 10'h1f0 == rs2[9:0] ? coeffs_496 : _GEN_1495;
  wire [31:0] _GEN_1497 = 10'h1f1 == rs2[9:0] ? coeffs_497 : _GEN_1496;
  wire [31:0] _GEN_1498 = 10'h1f2 == rs2[9:0] ? coeffs_498 : _GEN_1497;
  wire [31:0] _GEN_1499 = 10'h1f3 == rs2[9:0] ? coeffs_499 : _GEN_1498;
  wire [31:0] _GEN_1500 = 10'h1f4 == rs2[9:0] ? coeffs_500 : _GEN_1499;
  wire [31:0] _GEN_1501 = 10'h1f5 == rs2[9:0] ? coeffs_501 : _GEN_1500;
  wire [31:0] _GEN_1502 = 10'h1f6 == rs2[9:0] ? coeffs_502 : _GEN_1501;
  wire [31:0] _GEN_1503 = 10'h1f7 == rs2[9:0] ? coeffs_503 : _GEN_1502;
  wire [31:0] _GEN_1504 = 10'h1f8 == rs2[9:0] ? coeffs_504 : _GEN_1503;
  wire [31:0] _GEN_1505 = 10'h1f9 == rs2[9:0] ? coeffs_505 : _GEN_1504;
  wire [31:0] _GEN_1506 = 10'h1fa == rs2[9:0] ? coeffs_506 : _GEN_1505;
  wire [31:0] _GEN_1507 = 10'h1fb == rs2[9:0] ? coeffs_507 : _GEN_1506;
  wire [31:0] _GEN_1508 = 10'h1fc == rs2[9:0] ? coeffs_508 : _GEN_1507;
  wire [31:0] _GEN_1509 = 10'h1fd == rs2[9:0] ? coeffs_509 : _GEN_1508;
  wire [31:0] _GEN_1510 = 10'h1fe == rs2[9:0] ? coeffs_510 : _GEN_1509;
  wire [31:0] _GEN_1511 = 10'h1ff == rs2[9:0] ? coeffs_511 : _GEN_1510;
  wire [31:0] _GEN_1512 = 10'h200 == rs2[9:0] ? coeffs_512 : _GEN_1511;
  wire [31:0] _GEN_1513 = 10'h201 == rs2[9:0] ? coeffs_513 : _GEN_1512;
  wire [31:0] _GEN_1514 = 10'h202 == rs2[9:0] ? coeffs_514 : _GEN_1513;
  wire [31:0] _GEN_1515 = 10'h203 == rs2[9:0] ? coeffs_515 : _GEN_1514;
  wire [31:0] _GEN_1516 = 10'h204 == rs2[9:0] ? coeffs_516 : _GEN_1515;
  wire [31:0] _GEN_1517 = 10'h205 == rs2[9:0] ? coeffs_517 : _GEN_1516;
  wire [31:0] _GEN_1518 = 10'h206 == rs2[9:0] ? coeffs_518 : _GEN_1517;
  wire [31:0] _GEN_1519 = 10'h207 == rs2[9:0] ? coeffs_519 : _GEN_1518;
  wire [31:0] _GEN_1520 = 10'h208 == rs2[9:0] ? coeffs_520 : _GEN_1519;
  wire [31:0] _GEN_1521 = 10'h209 == rs2[9:0] ? coeffs_521 : _GEN_1520;
  wire [31:0] _GEN_1522 = 10'h20a == rs2[9:0] ? coeffs_522 : _GEN_1521;
  wire [31:0] _GEN_1523 = 10'h20b == rs2[9:0] ? coeffs_523 : _GEN_1522;
  wire [31:0] _GEN_1524 = 10'h20c == rs2[9:0] ? coeffs_524 : _GEN_1523;
  wire [31:0] _GEN_1525 = 10'h20d == rs2[9:0] ? coeffs_525 : _GEN_1524;
  wire [31:0] _GEN_1526 = 10'h20e == rs2[9:0] ? coeffs_526 : _GEN_1525;
  wire [31:0] _GEN_1527 = 10'h20f == rs2[9:0] ? coeffs_527 : _GEN_1526;
  wire [31:0] _GEN_1528 = 10'h210 == rs2[9:0] ? coeffs_528 : _GEN_1527;
  wire [31:0] _GEN_1529 = 10'h211 == rs2[9:0] ? coeffs_529 : _GEN_1528;
  wire [31:0] _GEN_1530 = 10'h212 == rs2[9:0] ? coeffs_530 : _GEN_1529;
  wire [31:0] _GEN_1531 = 10'h213 == rs2[9:0] ? coeffs_531 : _GEN_1530;
  wire [31:0] _GEN_1532 = 10'h214 == rs2[9:0] ? coeffs_532 : _GEN_1531;
  wire [31:0] _GEN_1533 = 10'h215 == rs2[9:0] ? coeffs_533 : _GEN_1532;
  wire [31:0] _GEN_1534 = 10'h216 == rs2[9:0] ? coeffs_534 : _GEN_1533;
  wire [31:0] _GEN_1535 = 10'h217 == rs2[9:0] ? coeffs_535 : _GEN_1534;
  wire [31:0] _GEN_1536 = 10'h218 == rs2[9:0] ? coeffs_536 : _GEN_1535;
  wire [31:0] _GEN_1537 = 10'h219 == rs2[9:0] ? coeffs_537 : _GEN_1536;
  wire [31:0] _GEN_1538 = 10'h21a == rs2[9:0] ? coeffs_538 : _GEN_1537;
  wire [31:0] _GEN_1539 = 10'h21b == rs2[9:0] ? coeffs_539 : _GEN_1538;
  wire [31:0] _GEN_1540 = 10'h21c == rs2[9:0] ? coeffs_540 : _GEN_1539;
  wire [31:0] _GEN_1541 = 10'h21d == rs2[9:0] ? coeffs_541 : _GEN_1540;
  wire [31:0] _GEN_1542 = 10'h21e == rs2[9:0] ? coeffs_542 : _GEN_1541;
  wire [31:0] _GEN_1543 = 10'h21f == rs2[9:0] ? coeffs_543 : _GEN_1542;
  wire [31:0] _GEN_1544 = 10'h220 == rs2[9:0] ? coeffs_544 : _GEN_1543;
  wire [31:0] _GEN_1545 = 10'h221 == rs2[9:0] ? coeffs_545 : _GEN_1544;
  wire [31:0] _GEN_1546 = 10'h222 == rs2[9:0] ? coeffs_546 : _GEN_1545;
  wire [31:0] _GEN_1547 = 10'h223 == rs2[9:0] ? coeffs_547 : _GEN_1546;
  wire [31:0] _GEN_1548 = 10'h224 == rs2[9:0] ? coeffs_548 : _GEN_1547;
  wire [31:0] _GEN_1549 = 10'h225 == rs2[9:0] ? coeffs_549 : _GEN_1548;
  wire [31:0] _GEN_1550 = 10'h226 == rs2[9:0] ? coeffs_550 : _GEN_1549;
  wire [31:0] _GEN_1551 = 10'h227 == rs2[9:0] ? coeffs_551 : _GEN_1550;
  wire [31:0] _GEN_1552 = 10'h228 == rs2[9:0] ? coeffs_552 : _GEN_1551;
  wire [31:0] _GEN_1553 = 10'h229 == rs2[9:0] ? coeffs_553 : _GEN_1552;
  wire [31:0] _GEN_1554 = 10'h22a == rs2[9:0] ? coeffs_554 : _GEN_1553;
  wire [31:0] _GEN_1555 = 10'h22b == rs2[9:0] ? coeffs_555 : _GEN_1554;
  wire [31:0] _GEN_1556 = 10'h22c == rs2[9:0] ? coeffs_556 : _GEN_1555;
  wire [31:0] _GEN_1557 = 10'h22d == rs2[9:0] ? coeffs_557 : _GEN_1556;
  wire [31:0] _GEN_1558 = 10'h22e == rs2[9:0] ? coeffs_558 : _GEN_1557;
  wire [31:0] _GEN_1559 = 10'h22f == rs2[9:0] ? coeffs_559 : _GEN_1558;
  wire [31:0] _GEN_1560 = 10'h230 == rs2[9:0] ? coeffs_560 : _GEN_1559;
  wire [31:0] _GEN_1561 = 10'h231 == rs2[9:0] ? coeffs_561 : _GEN_1560;
  wire [31:0] _GEN_1562 = 10'h232 == rs2[9:0] ? coeffs_562 : _GEN_1561;
  wire [31:0] _GEN_1563 = 10'h233 == rs2[9:0] ? coeffs_563 : _GEN_1562;
  wire [31:0] _GEN_1564 = 10'h234 == rs2[9:0] ? coeffs_564 : _GEN_1563;
  wire [31:0] _GEN_1565 = 10'h235 == rs2[9:0] ? coeffs_565 : _GEN_1564;
  wire [31:0] _GEN_1566 = 10'h236 == rs2[9:0] ? coeffs_566 : _GEN_1565;
  wire [31:0] _GEN_1567 = 10'h237 == rs2[9:0] ? coeffs_567 : _GEN_1566;
  wire [31:0] _GEN_1568 = 10'h238 == rs2[9:0] ? coeffs_568 : _GEN_1567;
  wire [31:0] _GEN_1569 = 10'h239 == rs2[9:0] ? coeffs_569 : _GEN_1568;
  wire [31:0] _GEN_1570 = 10'h23a == rs2[9:0] ? coeffs_570 : _GEN_1569;
  wire [31:0] _GEN_1571 = 10'h23b == rs2[9:0] ? coeffs_571 : _GEN_1570;
  wire [31:0] _GEN_1572 = 10'h23c == rs2[9:0] ? coeffs_572 : _GEN_1571;
  wire [31:0] _GEN_1573 = 10'h23d == rs2[9:0] ? coeffs_573 : _GEN_1572;
  wire [31:0] _GEN_1574 = 10'h23e == rs2[9:0] ? coeffs_574 : _GEN_1573;
  wire [31:0] _GEN_1575 = 10'h23f == rs2[9:0] ? coeffs_575 : _GEN_1574;
  wire [31:0] _GEN_1576 = 10'h240 == rs2[9:0] ? coeffs_576 : _GEN_1575;
  wire [31:0] _GEN_1577 = 10'h241 == rs2[9:0] ? coeffs_577 : _GEN_1576;
  wire [31:0] _GEN_1578 = 10'h242 == rs2[9:0] ? coeffs_578 : _GEN_1577;
  wire [31:0] _GEN_1579 = 10'h243 == rs2[9:0] ? coeffs_579 : _GEN_1578;
  wire [31:0] _GEN_1580 = 10'h244 == rs2[9:0] ? coeffs_580 : _GEN_1579;
  wire [31:0] _GEN_1581 = 10'h245 == rs2[9:0] ? coeffs_581 : _GEN_1580;
  wire [31:0] _GEN_1582 = 10'h246 == rs2[9:0] ? coeffs_582 : _GEN_1581;
  wire [31:0] _GEN_1583 = 10'h247 == rs2[9:0] ? coeffs_583 : _GEN_1582;
  wire [31:0] _GEN_1584 = 10'h248 == rs2[9:0] ? coeffs_584 : _GEN_1583;
  wire [31:0] _GEN_1585 = 10'h249 == rs2[9:0] ? coeffs_585 : _GEN_1584;
  wire [31:0] _GEN_1586 = 10'h24a == rs2[9:0] ? coeffs_586 : _GEN_1585;
  wire [31:0] _GEN_1587 = 10'h24b == rs2[9:0] ? coeffs_587 : _GEN_1586;
  wire [31:0] _GEN_1588 = 10'h24c == rs2[9:0] ? coeffs_588 : _GEN_1587;
  wire [31:0] _GEN_1589 = 10'h24d == rs2[9:0] ? coeffs_589 : _GEN_1588;
  wire [31:0] _GEN_1590 = 10'h24e == rs2[9:0] ? coeffs_590 : _GEN_1589;
  wire [31:0] _GEN_1591 = 10'h24f == rs2[9:0] ? coeffs_591 : _GEN_1590;
  wire [31:0] _GEN_1592 = 10'h250 == rs2[9:0] ? coeffs_592 : _GEN_1591;
  wire [31:0] _GEN_1593 = 10'h251 == rs2[9:0] ? coeffs_593 : _GEN_1592;
  wire [31:0] _GEN_1594 = 10'h252 == rs2[9:0] ? coeffs_594 : _GEN_1593;
  wire [31:0] _GEN_1595 = 10'h253 == rs2[9:0] ? coeffs_595 : _GEN_1594;
  wire [31:0] _GEN_1596 = 10'h254 == rs2[9:0] ? coeffs_596 : _GEN_1595;
  wire [31:0] _GEN_1597 = 10'h255 == rs2[9:0] ? coeffs_597 : _GEN_1596;
  wire [31:0] _GEN_1598 = 10'h256 == rs2[9:0] ? coeffs_598 : _GEN_1597;
  wire [31:0] _GEN_1599 = 10'h257 == rs2[9:0] ? coeffs_599 : _GEN_1598;
  wire [31:0] _GEN_1600 = 10'h258 == rs2[9:0] ? coeffs_600 : _GEN_1599;
  wire [31:0] _GEN_1601 = 10'h259 == rs2[9:0] ? coeffs_601 : _GEN_1600;
  wire [31:0] _GEN_1602 = 10'h25a == rs2[9:0] ? coeffs_602 : _GEN_1601;
  wire [31:0] _GEN_1603 = 10'h25b == rs2[9:0] ? coeffs_603 : _GEN_1602;
  wire [31:0] _GEN_1604 = 10'h25c == rs2[9:0] ? coeffs_604 : _GEN_1603;
  wire [31:0] _GEN_1605 = 10'h25d == rs2[9:0] ? coeffs_605 : _GEN_1604;
  wire [31:0] _GEN_1606 = 10'h25e == rs2[9:0] ? coeffs_606 : _GEN_1605;
  wire [31:0] _GEN_1607 = 10'h25f == rs2[9:0] ? coeffs_607 : _GEN_1606;
  wire [31:0] _GEN_1608 = 10'h260 == rs2[9:0] ? coeffs_608 : _GEN_1607;
  wire [31:0] _GEN_1609 = 10'h261 == rs2[9:0] ? coeffs_609 : _GEN_1608;
  wire [31:0] _GEN_1610 = 10'h262 == rs2[9:0] ? coeffs_610 : _GEN_1609;
  wire [31:0] _GEN_1611 = 10'h263 == rs2[9:0] ? coeffs_611 : _GEN_1610;
  wire [31:0] _GEN_1612 = 10'h264 == rs2[9:0] ? coeffs_612 : _GEN_1611;
  wire [31:0] _GEN_1613 = 10'h265 == rs2[9:0] ? coeffs_613 : _GEN_1612;
  wire [31:0] _GEN_1614 = 10'h266 == rs2[9:0] ? coeffs_614 : _GEN_1613;
  wire [31:0] _GEN_1615 = 10'h267 == rs2[9:0] ? coeffs_615 : _GEN_1614;
  wire [31:0] _GEN_1616 = 10'h268 == rs2[9:0] ? coeffs_616 : _GEN_1615;
  wire [31:0] _GEN_1617 = 10'h269 == rs2[9:0] ? coeffs_617 : _GEN_1616;
  wire [31:0] _GEN_1618 = 10'h26a == rs2[9:0] ? coeffs_618 : _GEN_1617;
  wire [31:0] _GEN_1619 = 10'h26b == rs2[9:0] ? coeffs_619 : _GEN_1618;
  wire [31:0] _GEN_1620 = 10'h26c == rs2[9:0] ? coeffs_620 : _GEN_1619;
  wire [31:0] _GEN_1621 = 10'h26d == rs2[9:0] ? coeffs_621 : _GEN_1620;
  wire [31:0] _GEN_1622 = 10'h26e == rs2[9:0] ? coeffs_622 : _GEN_1621;
  wire [31:0] _GEN_1623 = 10'h26f == rs2[9:0] ? coeffs_623 : _GEN_1622;
  wire [31:0] _GEN_1624 = 10'h270 == rs2[9:0] ? coeffs_624 : _GEN_1623;
  wire [31:0] _GEN_1625 = 10'h271 == rs2[9:0] ? coeffs_625 : _GEN_1624;
  wire [31:0] _GEN_1626 = 10'h272 == rs2[9:0] ? coeffs_626 : _GEN_1625;
  wire [31:0] _GEN_1627 = 10'h273 == rs2[9:0] ? coeffs_627 : _GEN_1626;
  wire [31:0] _GEN_1628 = 10'h274 == rs2[9:0] ? coeffs_628 : _GEN_1627;
  wire [31:0] _GEN_1629 = 10'h275 == rs2[9:0] ? coeffs_629 : _GEN_1628;
  wire [31:0] _GEN_1630 = 10'h276 == rs2[9:0] ? coeffs_630 : _GEN_1629;
  wire [31:0] _GEN_1631 = 10'h277 == rs2[9:0] ? coeffs_631 : _GEN_1630;
  wire [31:0] _GEN_1632 = 10'h278 == rs2[9:0] ? coeffs_632 : _GEN_1631;
  wire [31:0] _GEN_1633 = 10'h279 == rs2[9:0] ? coeffs_633 : _GEN_1632;
  wire [31:0] _GEN_1634 = 10'h27a == rs2[9:0] ? coeffs_634 : _GEN_1633;
  wire [31:0] _GEN_1635 = 10'h27b == rs2[9:0] ? coeffs_635 : _GEN_1634;
  wire [31:0] _GEN_1636 = 10'h27c == rs2[9:0] ? coeffs_636 : _GEN_1635;
  wire [31:0] _GEN_1637 = 10'h27d == rs2[9:0] ? coeffs_637 : _GEN_1636;
  wire [31:0] _GEN_1638 = 10'h27e == rs2[9:0] ? coeffs_638 : _GEN_1637;
  wire [31:0] _GEN_1639 = 10'h27f == rs2[9:0] ? coeffs_639 : _GEN_1638;
  wire [31:0] _GEN_1640 = 10'h280 == rs2[9:0] ? coeffs_640 : _GEN_1639;
  wire [31:0] _GEN_1641 = 10'h281 == rs2[9:0] ? coeffs_641 : _GEN_1640;
  wire [31:0] _GEN_1642 = 10'h282 == rs2[9:0] ? coeffs_642 : _GEN_1641;
  wire [31:0] _GEN_1643 = 10'h283 == rs2[9:0] ? coeffs_643 : _GEN_1642;
  wire [31:0] _GEN_1644 = 10'h284 == rs2[9:0] ? coeffs_644 : _GEN_1643;
  wire [31:0] _GEN_1645 = 10'h285 == rs2[9:0] ? coeffs_645 : _GEN_1644;
  wire [31:0] _GEN_1646 = 10'h286 == rs2[9:0] ? coeffs_646 : _GEN_1645;
  wire [31:0] _GEN_1647 = 10'h287 == rs2[9:0] ? coeffs_647 : _GEN_1646;
  wire [31:0] _GEN_1648 = 10'h288 == rs2[9:0] ? coeffs_648 : _GEN_1647;
  wire [31:0] _GEN_1649 = 10'h289 == rs2[9:0] ? coeffs_649 : _GEN_1648;
  wire [31:0] _GEN_1650 = 10'h28a == rs2[9:0] ? coeffs_650 : _GEN_1649;
  wire [31:0] _GEN_1651 = 10'h28b == rs2[9:0] ? coeffs_651 : _GEN_1650;
  wire [31:0] _GEN_1652 = 10'h28c == rs2[9:0] ? coeffs_652 : _GEN_1651;
  wire [31:0] _GEN_1653 = 10'h28d == rs2[9:0] ? coeffs_653 : _GEN_1652;
  wire [31:0] _GEN_1654 = 10'h28e == rs2[9:0] ? coeffs_654 : _GEN_1653;
  wire [31:0] _GEN_1655 = 10'h28f == rs2[9:0] ? coeffs_655 : _GEN_1654;
  wire [31:0] _GEN_1656 = 10'h290 == rs2[9:0] ? coeffs_656 : _GEN_1655;
  wire [31:0] _GEN_1657 = 10'h291 == rs2[9:0] ? coeffs_657 : _GEN_1656;
  wire [31:0] _GEN_1658 = 10'h292 == rs2[9:0] ? coeffs_658 : _GEN_1657;
  wire [31:0] _GEN_1659 = 10'h293 == rs2[9:0] ? coeffs_659 : _GEN_1658;
  wire [31:0] _GEN_1660 = 10'h294 == rs2[9:0] ? coeffs_660 : _GEN_1659;
  wire [31:0] _GEN_1661 = 10'h295 == rs2[9:0] ? coeffs_661 : _GEN_1660;
  wire [31:0] _GEN_1662 = 10'h296 == rs2[9:0] ? coeffs_662 : _GEN_1661;
  wire [31:0] _GEN_1663 = 10'h297 == rs2[9:0] ? coeffs_663 : _GEN_1662;
  wire [31:0] _GEN_1664 = 10'h298 == rs2[9:0] ? coeffs_664 : _GEN_1663;
  wire [31:0] _GEN_1665 = 10'h299 == rs2[9:0] ? coeffs_665 : _GEN_1664;
  wire [31:0] _GEN_1666 = 10'h29a == rs2[9:0] ? coeffs_666 : _GEN_1665;
  wire [31:0] _GEN_1667 = 10'h29b == rs2[9:0] ? coeffs_667 : _GEN_1666;
  wire [31:0] _GEN_1668 = 10'h29c == rs2[9:0] ? coeffs_668 : _GEN_1667;
  wire [31:0] _GEN_1669 = 10'h29d == rs2[9:0] ? coeffs_669 : _GEN_1668;
  wire [31:0] _GEN_1670 = 10'h29e == rs2[9:0] ? coeffs_670 : _GEN_1669;
  wire [31:0] _GEN_1671 = 10'h29f == rs2[9:0] ? coeffs_671 : _GEN_1670;
  wire [31:0] _GEN_1672 = 10'h2a0 == rs2[9:0] ? coeffs_672 : _GEN_1671;
  wire [31:0] _GEN_1673 = 10'h2a1 == rs2[9:0] ? coeffs_673 : _GEN_1672;
  wire [31:0] _GEN_1674 = 10'h2a2 == rs2[9:0] ? coeffs_674 : _GEN_1673;
  wire [31:0] _GEN_1675 = 10'h2a3 == rs2[9:0] ? coeffs_675 : _GEN_1674;
  wire [31:0] _GEN_1676 = 10'h2a4 == rs2[9:0] ? coeffs_676 : _GEN_1675;
  wire [31:0] _GEN_1677 = 10'h2a5 == rs2[9:0] ? coeffs_677 : _GEN_1676;
  wire [31:0] _GEN_1678 = 10'h2a6 == rs2[9:0] ? coeffs_678 : _GEN_1677;
  wire [31:0] _GEN_1679 = 10'h2a7 == rs2[9:0] ? coeffs_679 : _GEN_1678;
  wire [31:0] _GEN_1680 = 10'h2a8 == rs2[9:0] ? coeffs_680 : _GEN_1679;
  wire [31:0] _GEN_1681 = 10'h2a9 == rs2[9:0] ? coeffs_681 : _GEN_1680;
  wire [31:0] _GEN_1682 = 10'h2aa == rs2[9:0] ? coeffs_682 : _GEN_1681;
  wire [31:0] _GEN_1683 = 10'h2ab == rs2[9:0] ? coeffs_683 : _GEN_1682;
  wire [31:0] _GEN_1684 = 10'h2ac == rs2[9:0] ? coeffs_684 : _GEN_1683;
  wire [31:0] _GEN_1685 = 10'h2ad == rs2[9:0] ? coeffs_685 : _GEN_1684;
  wire [31:0] _GEN_1686 = 10'h2ae == rs2[9:0] ? coeffs_686 : _GEN_1685;
  wire [31:0] _GEN_1687 = 10'h2af == rs2[9:0] ? coeffs_687 : _GEN_1686;
  wire [31:0] _GEN_1688 = 10'h2b0 == rs2[9:0] ? coeffs_688 : _GEN_1687;
  wire [31:0] _GEN_1689 = 10'h2b1 == rs2[9:0] ? coeffs_689 : _GEN_1688;
  wire [31:0] _GEN_1690 = 10'h2b2 == rs2[9:0] ? coeffs_690 : _GEN_1689;
  wire [31:0] _GEN_1691 = 10'h2b3 == rs2[9:0] ? coeffs_691 : _GEN_1690;
  wire [31:0] _GEN_1692 = 10'h2b4 == rs2[9:0] ? coeffs_692 : _GEN_1691;
  wire [31:0] _GEN_1693 = 10'h2b5 == rs2[9:0] ? coeffs_693 : _GEN_1692;
  wire [31:0] _GEN_1694 = 10'h2b6 == rs2[9:0] ? coeffs_694 : _GEN_1693;
  wire [31:0] _GEN_1695 = 10'h2b7 == rs2[9:0] ? coeffs_695 : _GEN_1694;
  wire [31:0] _GEN_1696 = 10'h2b8 == rs2[9:0] ? coeffs_696 : _GEN_1695;
  wire [31:0] _GEN_1697 = 10'h2b9 == rs2[9:0] ? coeffs_697 : _GEN_1696;
  wire [31:0] _GEN_1698 = 10'h2ba == rs2[9:0] ? coeffs_698 : _GEN_1697;
  wire [31:0] _GEN_1699 = 10'h2bb == rs2[9:0] ? coeffs_699 : _GEN_1698;
  wire [31:0] _GEN_1700 = 10'h2bc == rs2[9:0] ? coeffs_700 : _GEN_1699;
  wire [31:0] _GEN_1701 = 10'h2bd == rs2[9:0] ? coeffs_701 : _GEN_1700;
  wire [31:0] _GEN_1702 = 10'h2be == rs2[9:0] ? coeffs_702 : _GEN_1701;
  wire [31:0] _GEN_1703 = 10'h2bf == rs2[9:0] ? coeffs_703 : _GEN_1702;
  wire [31:0] _GEN_1704 = 10'h2c0 == rs2[9:0] ? coeffs_704 : _GEN_1703;
  wire [31:0] _GEN_1705 = 10'h2c1 == rs2[9:0] ? coeffs_705 : _GEN_1704;
  wire [31:0] _GEN_1706 = 10'h2c2 == rs2[9:0] ? coeffs_706 : _GEN_1705;
  wire [31:0] _GEN_1707 = 10'h2c3 == rs2[9:0] ? coeffs_707 : _GEN_1706;
  wire [31:0] _GEN_1708 = 10'h2c4 == rs2[9:0] ? coeffs_708 : _GEN_1707;
  wire [31:0] _GEN_1709 = 10'h2c5 == rs2[9:0] ? coeffs_709 : _GEN_1708;
  wire [31:0] _GEN_1710 = 10'h2c6 == rs2[9:0] ? coeffs_710 : _GEN_1709;
  wire [31:0] _GEN_1711 = 10'h2c7 == rs2[9:0] ? coeffs_711 : _GEN_1710;
  wire [31:0] _GEN_1712 = 10'h2c8 == rs2[9:0] ? coeffs_712 : _GEN_1711;
  wire [31:0] _GEN_1713 = 10'h2c9 == rs2[9:0] ? coeffs_713 : _GEN_1712;
  wire [31:0] _GEN_1714 = 10'h2ca == rs2[9:0] ? coeffs_714 : _GEN_1713;
  wire [31:0] _GEN_1715 = 10'h2cb == rs2[9:0] ? coeffs_715 : _GEN_1714;
  wire [31:0] _GEN_1716 = 10'h2cc == rs2[9:0] ? coeffs_716 : _GEN_1715;
  wire [31:0] _GEN_1717 = 10'h2cd == rs2[9:0] ? coeffs_717 : _GEN_1716;
  wire [31:0] _GEN_1718 = 10'h2ce == rs2[9:0] ? coeffs_718 : _GEN_1717;
  wire [31:0] _GEN_1719 = 10'h2cf == rs2[9:0] ? coeffs_719 : _GEN_1718;
  wire [31:0] _GEN_1720 = 10'h2d0 == rs2[9:0] ? coeffs_720 : _GEN_1719;
  wire [31:0] _GEN_1721 = 10'h2d1 == rs2[9:0] ? coeffs_721 : _GEN_1720;
  wire [31:0] _GEN_1722 = 10'h2d2 == rs2[9:0] ? coeffs_722 : _GEN_1721;
  wire [31:0] _GEN_1723 = 10'h2d3 == rs2[9:0] ? coeffs_723 : _GEN_1722;
  wire [31:0] _GEN_1724 = 10'h2d4 == rs2[9:0] ? coeffs_724 : _GEN_1723;
  wire [31:0] _GEN_1725 = 10'h2d5 == rs2[9:0] ? coeffs_725 : _GEN_1724;
  wire [31:0] _GEN_1726 = 10'h2d6 == rs2[9:0] ? coeffs_726 : _GEN_1725;
  wire [31:0] _GEN_1727 = 10'h2d7 == rs2[9:0] ? coeffs_727 : _GEN_1726;
  wire [31:0] _GEN_1728 = 10'h2d8 == rs2[9:0] ? coeffs_728 : _GEN_1727;
  wire [31:0] _GEN_1729 = 10'h2d9 == rs2[9:0] ? coeffs_729 : _GEN_1728;
  wire [31:0] _GEN_1730 = 10'h2da == rs2[9:0] ? coeffs_730 : _GEN_1729;
  wire [31:0] _GEN_1731 = 10'h2db == rs2[9:0] ? coeffs_731 : _GEN_1730;
  wire [31:0] _GEN_1732 = 10'h2dc == rs2[9:0] ? coeffs_732 : _GEN_1731;
  wire [31:0] _GEN_1733 = 10'h2dd == rs2[9:0] ? coeffs_733 : _GEN_1732;
  wire [31:0] _GEN_1734 = 10'h2de == rs2[9:0] ? coeffs_734 : _GEN_1733;
  wire [31:0] _GEN_1735 = 10'h2df == rs2[9:0] ? coeffs_735 : _GEN_1734;
  wire [31:0] _GEN_1736 = 10'h2e0 == rs2[9:0] ? coeffs_736 : _GEN_1735;
  wire [31:0] _GEN_1737 = 10'h2e1 == rs2[9:0] ? coeffs_737 : _GEN_1736;
  wire [31:0] _GEN_1738 = 10'h2e2 == rs2[9:0] ? coeffs_738 : _GEN_1737;
  wire [31:0] _GEN_1739 = 10'h2e3 == rs2[9:0] ? coeffs_739 : _GEN_1738;
  wire [31:0] _GEN_1740 = 10'h2e4 == rs2[9:0] ? coeffs_740 : _GEN_1739;
  wire [31:0] _GEN_1741 = 10'h2e5 == rs2[9:0] ? coeffs_741 : _GEN_1740;
  wire [31:0] _GEN_1742 = 10'h2e6 == rs2[9:0] ? coeffs_742 : _GEN_1741;
  wire [31:0] _GEN_1743 = 10'h2e7 == rs2[9:0] ? coeffs_743 : _GEN_1742;
  wire [31:0] _GEN_1744 = 10'h2e8 == rs2[9:0] ? coeffs_744 : _GEN_1743;
  wire [31:0] _GEN_1745 = 10'h2e9 == rs2[9:0] ? coeffs_745 : _GEN_1744;
  wire [31:0] _GEN_1746 = 10'h2ea == rs2[9:0] ? coeffs_746 : _GEN_1745;
  wire [31:0] _GEN_1747 = 10'h2eb == rs2[9:0] ? coeffs_747 : _GEN_1746;
  wire [31:0] _GEN_1748 = 10'h2ec == rs2[9:0] ? coeffs_748 : _GEN_1747;
  wire [31:0] _GEN_1749 = 10'h2ed == rs2[9:0] ? coeffs_749 : _GEN_1748;
  wire [31:0] _GEN_1750 = 10'h2ee == rs2[9:0] ? coeffs_750 : _GEN_1749;
  wire [31:0] _GEN_1751 = 10'h2ef == rs2[9:0] ? coeffs_751 : _GEN_1750;
  wire [31:0] _GEN_1752 = 10'h2f0 == rs2[9:0] ? coeffs_752 : _GEN_1751;
  wire [31:0] _GEN_1753 = 10'h2f1 == rs2[9:0] ? coeffs_753 : _GEN_1752;
  wire [31:0] _GEN_1754 = 10'h2f2 == rs2[9:0] ? coeffs_754 : _GEN_1753;
  wire [31:0] _GEN_1755 = 10'h2f3 == rs2[9:0] ? coeffs_755 : _GEN_1754;
  wire [31:0] _GEN_1756 = 10'h2f4 == rs2[9:0] ? coeffs_756 : _GEN_1755;
  wire [31:0] _GEN_1757 = 10'h2f5 == rs2[9:0] ? coeffs_757 : _GEN_1756;
  wire [31:0] _GEN_1758 = 10'h2f6 == rs2[9:0] ? coeffs_758 : _GEN_1757;
  wire [31:0] _GEN_1759 = 10'h2f7 == rs2[9:0] ? coeffs_759 : _GEN_1758;
  wire [31:0] _GEN_1760 = 10'h2f8 == rs2[9:0] ? coeffs_760 : _GEN_1759;
  wire [31:0] _GEN_1761 = 10'h2f9 == rs2[9:0] ? coeffs_761 : _GEN_1760;
  wire [31:0] _GEN_1762 = 10'h2fa == rs2[9:0] ? coeffs_762 : _GEN_1761;
  wire [31:0] _GEN_1763 = 10'h2fb == rs2[9:0] ? coeffs_763 : _GEN_1762;
  wire [31:0] _GEN_1764 = 10'h2fc == rs2[9:0] ? coeffs_764 : _GEN_1763;
  wire [31:0] _GEN_1765 = 10'h2fd == rs2[9:0] ? coeffs_765 : _GEN_1764;
  wire [31:0] _GEN_1766 = 10'h2fe == rs2[9:0] ? coeffs_766 : _GEN_1765;
  wire [31:0] _GEN_1767 = 10'h2ff == rs2[9:0] ? coeffs_767 : _GEN_1766;
  wire [31:0] _GEN_1768 = 10'h300 == rs2[9:0] ? coeffs_768 : _GEN_1767;
  wire [31:0] _GEN_1769 = 10'h301 == rs2[9:0] ? coeffs_769 : _GEN_1768;
  wire [31:0] _GEN_1770 = 10'h302 == rs2[9:0] ? coeffs_770 : _GEN_1769;
  wire [31:0] _GEN_1771 = 10'h303 == rs2[9:0] ? coeffs_771 : _GEN_1770;
  wire [31:0] _GEN_1772 = 10'h304 == rs2[9:0] ? coeffs_772 : _GEN_1771;
  wire [31:0] _GEN_1773 = 10'h305 == rs2[9:0] ? coeffs_773 : _GEN_1772;
  wire [31:0] _GEN_1774 = 10'h306 == rs2[9:0] ? coeffs_774 : _GEN_1773;
  wire [31:0] _GEN_1775 = 10'h307 == rs2[9:0] ? coeffs_775 : _GEN_1774;
  wire [31:0] _GEN_1776 = 10'h308 == rs2[9:0] ? coeffs_776 : _GEN_1775;
  wire [31:0] _GEN_1777 = 10'h309 == rs2[9:0] ? coeffs_777 : _GEN_1776;
  wire [31:0] _GEN_1778 = 10'h30a == rs2[9:0] ? coeffs_778 : _GEN_1777;
  wire [31:0] _GEN_1779 = 10'h30b == rs2[9:0] ? coeffs_779 : _GEN_1778;
  wire [31:0] _GEN_1780 = 10'h30c == rs2[9:0] ? coeffs_780 : _GEN_1779;
  wire [31:0] _GEN_1781 = 10'h30d == rs2[9:0] ? coeffs_781 : _GEN_1780;
  wire [31:0] _GEN_1782 = 10'h30e == rs2[9:0] ? coeffs_782 : _GEN_1781;
  wire [31:0] _GEN_1783 = 10'h30f == rs2[9:0] ? coeffs_783 : _GEN_1782;
  wire [31:0] _GEN_1784 = 10'h310 == rs2[9:0] ? coeffs_784 : _GEN_1783;
  wire [31:0] _GEN_1785 = 10'h311 == rs2[9:0] ? coeffs_785 : _GEN_1784;
  wire [31:0] _GEN_1786 = 10'h312 == rs2[9:0] ? coeffs_786 : _GEN_1785;
  wire [31:0] _GEN_1787 = 10'h313 == rs2[9:0] ? coeffs_787 : _GEN_1786;
  wire [31:0] _GEN_1788 = 10'h314 == rs2[9:0] ? coeffs_788 : _GEN_1787;
  wire [31:0] _GEN_1789 = 10'h315 == rs2[9:0] ? coeffs_789 : _GEN_1788;
  wire [31:0] _GEN_1790 = 10'h316 == rs2[9:0] ? coeffs_790 : _GEN_1789;
  wire [31:0] _GEN_1791 = 10'h317 == rs2[9:0] ? coeffs_791 : _GEN_1790;
  wire [31:0] _GEN_1792 = 10'h318 == rs2[9:0] ? coeffs_792 : _GEN_1791;
  wire [31:0] _GEN_1793 = 10'h319 == rs2[9:0] ? coeffs_793 : _GEN_1792;
  wire [31:0] _GEN_1794 = 10'h31a == rs2[9:0] ? coeffs_794 : _GEN_1793;
  wire [31:0] _GEN_1795 = 10'h31b == rs2[9:0] ? coeffs_795 : _GEN_1794;
  wire [31:0] _GEN_1796 = 10'h31c == rs2[9:0] ? coeffs_796 : _GEN_1795;
  wire [31:0] _GEN_1797 = 10'h31d == rs2[9:0] ? coeffs_797 : _GEN_1796;
  wire [31:0] _GEN_1798 = 10'h31e == rs2[9:0] ? coeffs_798 : _GEN_1797;
  wire [31:0] _GEN_1799 = 10'h31f == rs2[9:0] ? coeffs_799 : _GEN_1798;
  wire [31:0] _GEN_1800 = 10'h320 == rs2[9:0] ? coeffs_800 : _GEN_1799;
  wire [31:0] _GEN_1801 = 10'h321 == rs2[9:0] ? coeffs_801 : _GEN_1800;
  wire [31:0] _GEN_1802 = 10'h322 == rs2[9:0] ? coeffs_802 : _GEN_1801;
  wire [31:0] _GEN_1803 = 10'h323 == rs2[9:0] ? coeffs_803 : _GEN_1802;
  wire [31:0] _GEN_1804 = 10'h324 == rs2[9:0] ? coeffs_804 : _GEN_1803;
  wire [31:0] _GEN_1805 = 10'h325 == rs2[9:0] ? coeffs_805 : _GEN_1804;
  wire [31:0] _GEN_1806 = 10'h326 == rs2[9:0] ? coeffs_806 : _GEN_1805;
  wire [31:0] _GEN_1807 = 10'h327 == rs2[9:0] ? coeffs_807 : _GEN_1806;
  wire [31:0] _GEN_1808 = 10'h328 == rs2[9:0] ? coeffs_808 : _GEN_1807;
  wire [31:0] _GEN_1809 = 10'h329 == rs2[9:0] ? coeffs_809 : _GEN_1808;
  wire [31:0] _GEN_1810 = 10'h32a == rs2[9:0] ? coeffs_810 : _GEN_1809;
  wire [31:0] _GEN_1811 = 10'h32b == rs2[9:0] ? coeffs_811 : _GEN_1810;
  wire [31:0] _GEN_1812 = 10'h32c == rs2[9:0] ? coeffs_812 : _GEN_1811;
  wire [31:0] _GEN_1813 = 10'h32d == rs2[9:0] ? coeffs_813 : _GEN_1812;
  wire [31:0] _GEN_1814 = 10'h32e == rs2[9:0] ? coeffs_814 : _GEN_1813;
  wire [31:0] _GEN_1815 = 10'h32f == rs2[9:0] ? coeffs_815 : _GEN_1814;
  wire [31:0] _GEN_1816 = 10'h330 == rs2[9:0] ? coeffs_816 : _GEN_1815;
  wire [31:0] _GEN_1817 = 10'h331 == rs2[9:0] ? coeffs_817 : _GEN_1816;
  wire [31:0] _GEN_1818 = 10'h332 == rs2[9:0] ? coeffs_818 : _GEN_1817;
  wire [31:0] _GEN_1819 = 10'h333 == rs2[9:0] ? coeffs_819 : _GEN_1818;
  wire [31:0] _GEN_1820 = 10'h334 == rs2[9:0] ? coeffs_820 : _GEN_1819;
  wire [31:0] _GEN_1821 = 10'h335 == rs2[9:0] ? coeffs_821 : _GEN_1820;
  wire [31:0] _GEN_1822 = 10'h336 == rs2[9:0] ? coeffs_822 : _GEN_1821;
  wire [31:0] _GEN_1823 = 10'h337 == rs2[9:0] ? coeffs_823 : _GEN_1822;
  wire [31:0] _GEN_1824 = 10'h338 == rs2[9:0] ? coeffs_824 : _GEN_1823;
  wire [31:0] _GEN_1825 = 10'h339 == rs2[9:0] ? coeffs_825 : _GEN_1824;
  wire [31:0] _GEN_1826 = 10'h33a == rs2[9:0] ? coeffs_826 : _GEN_1825;
  wire [31:0] _GEN_1827 = 10'h33b == rs2[9:0] ? coeffs_827 : _GEN_1826;
  wire [31:0] _GEN_1828 = 10'h33c == rs2[9:0] ? coeffs_828 : _GEN_1827;
  wire [31:0] _GEN_1829 = 10'h33d == rs2[9:0] ? coeffs_829 : _GEN_1828;
  wire [31:0] _GEN_1830 = 10'h33e == rs2[9:0] ? coeffs_830 : _GEN_1829;
  wire [31:0] _GEN_1831 = 10'h33f == rs2[9:0] ? coeffs_831 : _GEN_1830;
  wire [31:0] _GEN_1832 = 10'h340 == rs2[9:0] ? coeffs_832 : _GEN_1831;
  wire [31:0] _GEN_1833 = 10'h341 == rs2[9:0] ? coeffs_833 : _GEN_1832;
  wire [31:0] _GEN_1834 = 10'h342 == rs2[9:0] ? coeffs_834 : _GEN_1833;
  wire [31:0] _GEN_1835 = 10'h343 == rs2[9:0] ? coeffs_835 : _GEN_1834;
  wire [31:0] _GEN_1836 = 10'h344 == rs2[9:0] ? coeffs_836 : _GEN_1835;
  wire [31:0] _GEN_1837 = 10'h345 == rs2[9:0] ? coeffs_837 : _GEN_1836;
  wire [31:0] _GEN_1838 = 10'h346 == rs2[9:0] ? coeffs_838 : _GEN_1837;
  wire [31:0] _GEN_1839 = 10'h347 == rs2[9:0] ? coeffs_839 : _GEN_1838;
  wire [31:0] _GEN_1840 = 10'h348 == rs2[9:0] ? coeffs_840 : _GEN_1839;
  wire [31:0] _GEN_1841 = 10'h349 == rs2[9:0] ? coeffs_841 : _GEN_1840;
  wire [31:0] _GEN_1842 = 10'h34a == rs2[9:0] ? coeffs_842 : _GEN_1841;
  wire [31:0] _GEN_1843 = 10'h34b == rs2[9:0] ? coeffs_843 : _GEN_1842;
  wire [31:0] _GEN_1844 = 10'h34c == rs2[9:0] ? coeffs_844 : _GEN_1843;
  wire [31:0] _GEN_1845 = 10'h34d == rs2[9:0] ? coeffs_845 : _GEN_1844;
  wire [31:0] _GEN_1846 = 10'h34e == rs2[9:0] ? coeffs_846 : _GEN_1845;
  wire [31:0] _GEN_1847 = 10'h34f == rs2[9:0] ? coeffs_847 : _GEN_1846;
  wire [31:0] _GEN_1848 = 10'h350 == rs2[9:0] ? coeffs_848 : _GEN_1847;
  wire [31:0] _GEN_1849 = 10'h351 == rs2[9:0] ? coeffs_849 : _GEN_1848;
  wire [31:0] _GEN_1850 = 10'h352 == rs2[9:0] ? coeffs_850 : _GEN_1849;
  wire [31:0] _GEN_1851 = 10'h353 == rs2[9:0] ? coeffs_851 : _GEN_1850;
  wire [31:0] _GEN_1852 = 10'h354 == rs2[9:0] ? coeffs_852 : _GEN_1851;
  wire [31:0] _GEN_1853 = 10'h355 == rs2[9:0] ? coeffs_853 : _GEN_1852;
  wire [31:0] _GEN_1854 = 10'h356 == rs2[9:0] ? coeffs_854 : _GEN_1853;
  wire [31:0] _GEN_1855 = 10'h357 == rs2[9:0] ? coeffs_855 : _GEN_1854;
  wire [31:0] _GEN_1856 = 10'h358 == rs2[9:0] ? coeffs_856 : _GEN_1855;
  wire [31:0] _GEN_1857 = 10'h359 == rs2[9:0] ? coeffs_857 : _GEN_1856;
  wire [31:0] _GEN_1858 = 10'h35a == rs2[9:0] ? coeffs_858 : _GEN_1857;
  wire [31:0] _GEN_1859 = 10'h35b == rs2[9:0] ? coeffs_859 : _GEN_1858;
  wire [31:0] _GEN_1860 = 10'h35c == rs2[9:0] ? coeffs_860 : _GEN_1859;
  wire [31:0] _GEN_1861 = 10'h35d == rs2[9:0] ? coeffs_861 : _GEN_1860;
  wire [31:0] _GEN_1862 = 10'h35e == rs2[9:0] ? coeffs_862 : _GEN_1861;
  wire [31:0] _GEN_1863 = 10'h35f == rs2[9:0] ? coeffs_863 : _GEN_1862;
  wire [31:0] _GEN_1864 = 10'h360 == rs2[9:0] ? coeffs_864 : _GEN_1863;
  wire [31:0] _GEN_1865 = 10'h361 == rs2[9:0] ? coeffs_865 : _GEN_1864;
  wire [31:0] _GEN_1866 = 10'h362 == rs2[9:0] ? coeffs_866 : _GEN_1865;
  wire [31:0] _GEN_1867 = 10'h363 == rs2[9:0] ? coeffs_867 : _GEN_1866;
  wire [31:0] _GEN_1868 = 10'h364 == rs2[9:0] ? coeffs_868 : _GEN_1867;
  wire [31:0] _GEN_1869 = 10'h365 == rs2[9:0] ? coeffs_869 : _GEN_1868;
  wire [31:0] _GEN_1870 = 10'h366 == rs2[9:0] ? coeffs_870 : _GEN_1869;
  wire [31:0] _GEN_1871 = 10'h367 == rs2[9:0] ? coeffs_871 : _GEN_1870;
  wire [31:0] _GEN_1872 = 10'h368 == rs2[9:0] ? coeffs_872 : _GEN_1871;
  wire [31:0] _GEN_1873 = 10'h369 == rs2[9:0] ? coeffs_873 : _GEN_1872;
  wire [31:0] _GEN_1874 = 10'h36a == rs2[9:0] ? coeffs_874 : _GEN_1873;
  wire [31:0] _GEN_1875 = 10'h36b == rs2[9:0] ? coeffs_875 : _GEN_1874;
  wire [31:0] _GEN_1876 = 10'h36c == rs2[9:0] ? coeffs_876 : _GEN_1875;
  wire [31:0] _GEN_1877 = 10'h36d == rs2[9:0] ? coeffs_877 : _GEN_1876;
  wire [31:0] _GEN_1878 = 10'h36e == rs2[9:0] ? coeffs_878 : _GEN_1877;
  wire [31:0] _GEN_1879 = 10'h36f == rs2[9:0] ? coeffs_879 : _GEN_1878;
  wire [31:0] _GEN_1880 = 10'h370 == rs2[9:0] ? coeffs_880 : _GEN_1879;
  wire [31:0] _GEN_1881 = 10'h371 == rs2[9:0] ? coeffs_881 : _GEN_1880;
  wire [31:0] _GEN_1882 = 10'h372 == rs2[9:0] ? coeffs_882 : _GEN_1881;
  wire [31:0] _GEN_1883 = 10'h373 == rs2[9:0] ? coeffs_883 : _GEN_1882;
  wire [31:0] _GEN_1884 = 10'h374 == rs2[9:0] ? coeffs_884 : _GEN_1883;
  wire [31:0] _GEN_1885 = 10'h375 == rs2[9:0] ? coeffs_885 : _GEN_1884;
  wire [31:0] _GEN_1886 = 10'h376 == rs2[9:0] ? coeffs_886 : _GEN_1885;
  wire [31:0] _GEN_1887 = 10'h377 == rs2[9:0] ? coeffs_887 : _GEN_1886;
  wire [31:0] _GEN_1888 = 10'h378 == rs2[9:0] ? coeffs_888 : _GEN_1887;
  wire [31:0] _GEN_1889 = 10'h379 == rs2[9:0] ? coeffs_889 : _GEN_1888;
  wire [31:0] _GEN_1890 = 10'h37a == rs2[9:0] ? coeffs_890 : _GEN_1889;
  wire [31:0] _GEN_1891 = 10'h37b == rs2[9:0] ? coeffs_891 : _GEN_1890;
  wire [31:0] _GEN_1892 = 10'h37c == rs2[9:0] ? coeffs_892 : _GEN_1891;
  wire [31:0] _GEN_1893 = 10'h37d == rs2[9:0] ? coeffs_893 : _GEN_1892;
  wire [31:0] _GEN_1894 = 10'h37e == rs2[9:0] ? coeffs_894 : _GEN_1893;
  wire [31:0] _GEN_1895 = 10'h37f == rs2[9:0] ? coeffs_895 : _GEN_1894;
  wire [31:0] _GEN_1896 = 10'h380 == rs2[9:0] ? coeffs_896 : _GEN_1895;
  wire [31:0] _GEN_1897 = 10'h381 == rs2[9:0] ? coeffs_897 : _GEN_1896;
  wire [31:0] _GEN_1898 = 10'h382 == rs2[9:0] ? coeffs_898 : _GEN_1897;
  wire [31:0] _GEN_1899 = 10'h383 == rs2[9:0] ? coeffs_899 : _GEN_1898;
  wire [31:0] _GEN_1900 = 10'h384 == rs2[9:0] ? coeffs_900 : _GEN_1899;
  wire [31:0] _GEN_1901 = 10'h385 == rs2[9:0] ? coeffs_901 : _GEN_1900;
  wire [31:0] _GEN_1902 = 10'h386 == rs2[9:0] ? coeffs_902 : _GEN_1901;
  wire [31:0] _GEN_1903 = 10'h387 == rs2[9:0] ? coeffs_903 : _GEN_1902;
  wire [31:0] _GEN_1904 = 10'h388 == rs2[9:0] ? coeffs_904 : _GEN_1903;
  wire [31:0] _GEN_1905 = 10'h389 == rs2[9:0] ? coeffs_905 : _GEN_1904;
  wire [31:0] _GEN_1906 = 10'h38a == rs2[9:0] ? coeffs_906 : _GEN_1905;
  wire [31:0] _GEN_1907 = 10'h38b == rs2[9:0] ? coeffs_907 : _GEN_1906;
  wire [31:0] _GEN_1908 = 10'h38c == rs2[9:0] ? coeffs_908 : _GEN_1907;
  wire [31:0] _GEN_1909 = 10'h38d == rs2[9:0] ? coeffs_909 : _GEN_1908;
  wire [31:0] _GEN_1910 = 10'h38e == rs2[9:0] ? coeffs_910 : _GEN_1909;
  wire [31:0] _GEN_1911 = 10'h38f == rs2[9:0] ? coeffs_911 : _GEN_1910;
  wire [31:0] _GEN_1912 = 10'h390 == rs2[9:0] ? coeffs_912 : _GEN_1911;
  wire [31:0] _GEN_1913 = 10'h391 == rs2[9:0] ? coeffs_913 : _GEN_1912;
  wire [31:0] _GEN_1914 = 10'h392 == rs2[9:0] ? coeffs_914 : _GEN_1913;
  wire [31:0] _GEN_1915 = 10'h393 == rs2[9:0] ? coeffs_915 : _GEN_1914;
  wire [31:0] _GEN_1916 = 10'h394 == rs2[9:0] ? coeffs_916 : _GEN_1915;
  wire [31:0] _GEN_1917 = 10'h395 == rs2[9:0] ? coeffs_917 : _GEN_1916;
  wire [31:0] _GEN_1918 = 10'h396 == rs2[9:0] ? coeffs_918 : _GEN_1917;
  wire [31:0] _GEN_1919 = 10'h397 == rs2[9:0] ? coeffs_919 : _GEN_1918;
  wire [31:0] _GEN_1920 = 10'h398 == rs2[9:0] ? coeffs_920 : _GEN_1919;
  wire [31:0] _GEN_1921 = 10'h399 == rs2[9:0] ? coeffs_921 : _GEN_1920;
  wire [31:0] _GEN_1922 = 10'h39a == rs2[9:0] ? coeffs_922 : _GEN_1921;
  wire [31:0] _GEN_1923 = 10'h39b == rs2[9:0] ? coeffs_923 : _GEN_1922;
  wire [31:0] _GEN_1924 = 10'h39c == rs2[9:0] ? coeffs_924 : _GEN_1923;
  wire [31:0] _GEN_1925 = 10'h39d == rs2[9:0] ? coeffs_925 : _GEN_1924;
  wire [31:0] _GEN_1926 = 10'h39e == rs2[9:0] ? coeffs_926 : _GEN_1925;
  wire [31:0] _GEN_1927 = 10'h39f == rs2[9:0] ? coeffs_927 : _GEN_1926;
  wire [31:0] _GEN_1928 = 10'h3a0 == rs2[9:0] ? coeffs_928 : _GEN_1927;
  wire [31:0] _GEN_1929 = 10'h3a1 == rs2[9:0] ? coeffs_929 : _GEN_1928;
  wire [31:0] _GEN_1930 = 10'h3a2 == rs2[9:0] ? coeffs_930 : _GEN_1929;
  wire [31:0] _GEN_1931 = 10'h3a3 == rs2[9:0] ? coeffs_931 : _GEN_1930;
  wire [31:0] _GEN_1932 = 10'h3a4 == rs2[9:0] ? coeffs_932 : _GEN_1931;
  wire [31:0] _GEN_1933 = 10'h3a5 == rs2[9:0] ? coeffs_933 : _GEN_1932;
  wire [31:0] _GEN_1934 = 10'h3a6 == rs2[9:0] ? coeffs_934 : _GEN_1933;
  wire [31:0] _GEN_1935 = 10'h3a7 == rs2[9:0] ? coeffs_935 : _GEN_1934;
  wire [31:0] _GEN_1936 = 10'h3a8 == rs2[9:0] ? coeffs_936 : _GEN_1935;
  wire [31:0] _GEN_1937 = 10'h3a9 == rs2[9:0] ? coeffs_937 : _GEN_1936;
  wire [31:0] _GEN_1938 = 10'h3aa == rs2[9:0] ? coeffs_938 : _GEN_1937;
  wire [31:0] _GEN_1939 = 10'h3ab == rs2[9:0] ? coeffs_939 : _GEN_1938;
  wire [31:0] _GEN_1940 = 10'h3ac == rs2[9:0] ? coeffs_940 : _GEN_1939;
  wire [31:0] _GEN_1941 = 10'h3ad == rs2[9:0] ? coeffs_941 : _GEN_1940;
  wire [31:0] _GEN_1942 = 10'h3ae == rs2[9:0] ? coeffs_942 : _GEN_1941;
  wire [31:0] _GEN_1943 = 10'h3af == rs2[9:0] ? coeffs_943 : _GEN_1942;
  wire [31:0] _GEN_1944 = 10'h3b0 == rs2[9:0] ? coeffs_944 : _GEN_1943;
  wire [31:0] _GEN_1945 = 10'h3b1 == rs2[9:0] ? coeffs_945 : _GEN_1944;
  wire [31:0] _GEN_1946 = 10'h3b2 == rs2[9:0] ? coeffs_946 : _GEN_1945;
  wire [31:0] _GEN_1947 = 10'h3b3 == rs2[9:0] ? coeffs_947 : _GEN_1946;
  wire [31:0] _GEN_1948 = 10'h3b4 == rs2[9:0] ? coeffs_948 : _GEN_1947;
  wire [31:0] _GEN_1949 = 10'h3b5 == rs2[9:0] ? coeffs_949 : _GEN_1948;
  wire [31:0] _GEN_1950 = 10'h3b6 == rs2[9:0] ? coeffs_950 : _GEN_1949;
  wire [31:0] _GEN_1951 = 10'h3b7 == rs2[9:0] ? coeffs_951 : _GEN_1950;
  wire [31:0] _GEN_1952 = 10'h3b8 == rs2[9:0] ? coeffs_952 : _GEN_1951;
  wire [31:0] _GEN_1953 = 10'h3b9 == rs2[9:0] ? coeffs_953 : _GEN_1952;
  wire [31:0] _GEN_1954 = 10'h3ba == rs2[9:0] ? coeffs_954 : _GEN_1953;
  wire [31:0] _GEN_1955 = 10'h3bb == rs2[9:0] ? coeffs_955 : _GEN_1954;
  wire [31:0] _GEN_1956 = 10'h3bc == rs2[9:0] ? coeffs_956 : _GEN_1955;
  wire [31:0] _GEN_1957 = 10'h3bd == rs2[9:0] ? coeffs_957 : _GEN_1956;
  wire [31:0] _GEN_1958 = 10'h3be == rs2[9:0] ? coeffs_958 : _GEN_1957;
  wire [31:0] _GEN_1959 = 10'h3bf == rs2[9:0] ? coeffs_959 : _GEN_1958;
  wire [31:0] _GEN_1960 = 10'h3c0 == rs2[9:0] ? coeffs_960 : _GEN_1959;
  wire [31:0] _GEN_1961 = 10'h3c1 == rs2[9:0] ? coeffs_961 : _GEN_1960;
  wire [31:0] _GEN_1962 = 10'h3c2 == rs2[9:0] ? coeffs_962 : _GEN_1961;
  wire [31:0] _GEN_1963 = 10'h3c3 == rs2[9:0] ? coeffs_963 : _GEN_1962;
  wire [31:0] _GEN_1964 = 10'h3c4 == rs2[9:0] ? coeffs_964 : _GEN_1963;
  wire [31:0] _GEN_1965 = 10'h3c5 == rs2[9:0] ? coeffs_965 : _GEN_1964;
  wire [31:0] _GEN_1966 = 10'h3c6 == rs2[9:0] ? coeffs_966 : _GEN_1965;
  wire [31:0] _GEN_1967 = 10'h3c7 == rs2[9:0] ? coeffs_967 : _GEN_1966;
  wire [31:0] _GEN_1968 = 10'h3c8 == rs2[9:0] ? coeffs_968 : _GEN_1967;
  wire [31:0] _GEN_1969 = 10'h3c9 == rs2[9:0] ? coeffs_969 : _GEN_1968;
  wire [31:0] _GEN_1970 = 10'h3ca == rs2[9:0] ? coeffs_970 : _GEN_1969;
  wire [31:0] _GEN_1971 = 10'h3cb == rs2[9:0] ? coeffs_971 : _GEN_1970;
  wire [31:0] _GEN_1972 = 10'h3cc == rs2[9:0] ? coeffs_972 : _GEN_1971;
  wire [31:0] _GEN_1973 = 10'h3cd == rs2[9:0] ? coeffs_973 : _GEN_1972;
  wire [31:0] _GEN_1974 = 10'h3ce == rs2[9:0] ? coeffs_974 : _GEN_1973;
  wire [31:0] _GEN_1975 = 10'h3cf == rs2[9:0] ? coeffs_975 : _GEN_1974;
  wire [31:0] _GEN_1976 = 10'h3d0 == rs2[9:0] ? coeffs_976 : _GEN_1975;
  wire [31:0] _GEN_1977 = 10'h3d1 == rs2[9:0] ? coeffs_977 : _GEN_1976;
  wire [31:0] _GEN_1978 = 10'h3d2 == rs2[9:0] ? coeffs_978 : _GEN_1977;
  wire [31:0] _GEN_1979 = 10'h3d3 == rs2[9:0] ? coeffs_979 : _GEN_1978;
  wire [31:0] _GEN_1980 = 10'h3d4 == rs2[9:0] ? coeffs_980 : _GEN_1979;
  wire [31:0] _GEN_1981 = 10'h3d5 == rs2[9:0] ? coeffs_981 : _GEN_1980;
  wire [31:0] _GEN_1982 = 10'h3d6 == rs2[9:0] ? coeffs_982 : _GEN_1981;
  wire [31:0] _GEN_1983 = 10'h3d7 == rs2[9:0] ? coeffs_983 : _GEN_1982;
  wire [31:0] _GEN_1984 = 10'h3d8 == rs2[9:0] ? coeffs_984 : _GEN_1983;
  wire [31:0] _GEN_1985 = 10'h3d9 == rs2[9:0] ? coeffs_985 : _GEN_1984;
  wire [31:0] _GEN_1986 = 10'h3da == rs2[9:0] ? coeffs_986 : _GEN_1985;
  wire [31:0] _GEN_1987 = 10'h3db == rs2[9:0] ? coeffs_987 : _GEN_1986;
  wire [31:0] _GEN_1988 = 10'h3dc == rs2[9:0] ? coeffs_988 : _GEN_1987;
  wire [31:0] _GEN_1989 = 10'h3dd == rs2[9:0] ? coeffs_989 : _GEN_1988;
  wire [31:0] _GEN_1990 = 10'h3de == rs2[9:0] ? coeffs_990 : _GEN_1989;
  wire [31:0] _GEN_1991 = 10'h3df == rs2[9:0] ? coeffs_991 : _GEN_1990;
  wire [31:0] _GEN_1992 = 10'h3e0 == rs2[9:0] ? coeffs_992 : _GEN_1991;
  wire [31:0] _GEN_1993 = 10'h3e1 == rs2[9:0] ? coeffs_993 : _GEN_1992;
  wire [31:0] _GEN_1994 = 10'h3e2 == rs2[9:0] ? coeffs_994 : _GEN_1993;
  wire [31:0] _GEN_1995 = 10'h3e3 == rs2[9:0] ? coeffs_995 : _GEN_1994;
  wire [31:0] _GEN_1996 = 10'h3e4 == rs2[9:0] ? coeffs_996 : _GEN_1995;
  wire [31:0] _GEN_1997 = 10'h3e5 == rs2[9:0] ? coeffs_997 : _GEN_1996;
  wire [31:0] _GEN_1998 = 10'h3e6 == rs2[9:0] ? coeffs_998 : _GEN_1997;
  wire [31:0] _GEN_1999 = 10'h3e7 == rs2[9:0] ? coeffs_999 : _GEN_1998;
  wire [63:0] _result_T_1 = data_0 * coeffs_0;
  wire [63:0] _result_T_2 = data_1 * coeffs_1;
  wire [63:0] _result_T_3 = data_2 * coeffs_2;
  wire [63:0] _result_T_4 = data_3 * coeffs_3;
  wire [63:0] _result_T_5 = data_4 * coeffs_4;
  wire [63:0] _result_T_6 = data_5 * coeffs_5;
  wire [63:0] _result_T_7 = data_6 * coeffs_6;
  wire [63:0] _result_T_8 = data_7 * coeffs_7;
  wire [63:0] _result_T_9 = data_8 * coeffs_8;
  wire [63:0] _result_T_10 = data_9 * coeffs_9;
  wire [63:0] _result_T_11 = data_10 * coeffs_10;
  wire [63:0] _result_T_12 = data_11 * coeffs_11;
  wire [63:0] _result_T_13 = data_12 * coeffs_12;
  wire [63:0] _result_T_14 = data_13 * coeffs_13;
  wire [63:0] _result_T_15 = data_14 * coeffs_14;
  wire [63:0] _result_T_16 = data_15 * coeffs_15;
  wire [63:0] _result_T_17 = data_16 * coeffs_16;
  wire [63:0] _result_T_18 = data_17 * coeffs_17;
  wire [63:0] _result_T_19 = data_18 * coeffs_18;
  wire [63:0] _result_T_20 = data_19 * coeffs_19;
  wire [63:0] _result_T_21 = data_20 * coeffs_20;
  wire [63:0] _result_T_22 = data_21 * coeffs_21;
  wire [63:0] _result_T_23 = data_22 * coeffs_22;
  wire [63:0] _result_T_24 = data_23 * coeffs_23;
  wire [63:0] _result_T_25 = data_24 * coeffs_24;
  wire [63:0] _result_T_26 = data_25 * coeffs_25;
  wire [63:0] _result_T_27 = data_26 * coeffs_26;
  wire [63:0] _result_T_28 = data_27 * coeffs_27;
  wire [63:0] _result_T_29 = data_28 * coeffs_28;
  wire [63:0] _result_T_30 = data_29 * coeffs_29;
  wire [63:0] _result_T_31 = data_30 * coeffs_30;
  wire [63:0] _result_T_32 = data_31 * coeffs_31;
  wire [63:0] _result_T_33 = data_32 * coeffs_32;
  wire [63:0] _result_T_34 = data_33 * coeffs_33;
  wire [63:0] _result_T_35 = data_34 * coeffs_34;
  wire [63:0] _result_T_36 = data_35 * coeffs_35;
  wire [63:0] _result_T_37 = data_36 * coeffs_36;
  wire [63:0] _result_T_38 = data_37 * coeffs_37;
  wire [63:0] _result_T_39 = data_38 * coeffs_38;
  wire [63:0] _result_T_40 = data_39 * coeffs_39;
  wire [63:0] _result_T_41 = data_40 * coeffs_40;
  wire [63:0] _result_T_42 = data_41 * coeffs_41;
  wire [63:0] _result_T_43 = data_42 * coeffs_42;
  wire [63:0] _result_T_44 = data_43 * coeffs_43;
  wire [63:0] _result_T_45 = data_44 * coeffs_44;
  wire [63:0] _result_T_46 = data_45 * coeffs_45;
  wire [63:0] _result_T_47 = data_46 * coeffs_46;
  wire [63:0] _result_T_48 = data_47 * coeffs_47;
  wire [63:0] _result_T_49 = data_48 * coeffs_48;
  wire [63:0] _result_T_50 = data_49 * coeffs_49;
  wire [63:0] _result_T_51 = data_50 * coeffs_50;
  wire [63:0] _result_T_52 = data_51 * coeffs_51;
  wire [63:0] _result_T_53 = data_52 * coeffs_52;
  wire [63:0] _result_T_54 = data_53 * coeffs_53;
  wire [63:0] _result_T_55 = data_54 * coeffs_54;
  wire [63:0] _result_T_56 = data_55 * coeffs_55;
  wire [63:0] _result_T_57 = data_56 * coeffs_56;
  wire [63:0] _result_T_58 = data_57 * coeffs_57;
  wire [63:0] _result_T_59 = data_58 * coeffs_58;
  wire [63:0] _result_T_60 = data_59 * coeffs_59;
  wire [63:0] _result_T_61 = data_60 * coeffs_60;
  wire [63:0] _result_T_62 = data_61 * coeffs_61;
  wire [63:0] _result_T_63 = data_62 * coeffs_62;
  wire [63:0] _result_T_64 = data_63 * coeffs_63;
  wire [63:0] _result_T_65 = data_64 * coeffs_64;
  wire [63:0] _result_T_66 = data_65 * coeffs_65;
  wire [63:0] _result_T_67 = data_66 * coeffs_66;
  wire [63:0] _result_T_68 = data_67 * coeffs_67;
  wire [63:0] _result_T_69 = data_68 * coeffs_68;
  wire [63:0] _result_T_70 = data_69 * coeffs_69;
  wire [63:0] _result_T_71 = data_70 * coeffs_70;
  wire [63:0] _result_T_72 = data_71 * coeffs_71;
  wire [63:0] _result_T_73 = data_72 * coeffs_72;
  wire [63:0] _result_T_74 = data_73 * coeffs_73;
  wire [63:0] _result_T_75 = data_74 * coeffs_74;
  wire [63:0] _result_T_76 = data_75 * coeffs_75;
  wire [63:0] _result_T_77 = data_76 * coeffs_76;
  wire [63:0] _result_T_78 = data_77 * coeffs_77;
  wire [63:0] _result_T_79 = data_78 * coeffs_78;
  wire [63:0] _result_T_80 = data_79 * coeffs_79;
  wire [63:0] _result_T_81 = data_80 * coeffs_80;
  wire [63:0] _result_T_82 = data_81 * coeffs_81;
  wire [63:0] _result_T_83 = data_82 * coeffs_82;
  wire [63:0] _result_T_84 = data_83 * coeffs_83;
  wire [63:0] _result_T_85 = data_84 * coeffs_84;
  wire [63:0] _result_T_86 = data_85 * coeffs_85;
  wire [63:0] _result_T_87 = data_86 * coeffs_86;
  wire [63:0] _result_T_88 = data_87 * coeffs_87;
  wire [63:0] _result_T_89 = data_88 * coeffs_88;
  wire [63:0] _result_T_90 = data_89 * coeffs_89;
  wire [63:0] _result_T_91 = data_90 * coeffs_90;
  wire [63:0] _result_T_92 = data_91 * coeffs_91;
  wire [63:0] _result_T_93 = data_92 * coeffs_92;
  wire [63:0] _result_T_94 = data_93 * coeffs_93;
  wire [63:0] _result_T_95 = data_94 * coeffs_94;
  wire [63:0] _result_T_96 = data_95 * coeffs_95;
  wire [63:0] _result_T_97 = data_96 * coeffs_96;
  wire [63:0] _result_T_98 = data_97 * coeffs_97;
  wire [63:0] _result_T_99 = data_98 * coeffs_98;
  wire [63:0] _result_T_100 = data_99 * coeffs_99;
  wire [63:0] _result_T_101 = data_100 * coeffs_100;
  wire [63:0] _result_T_102 = data_101 * coeffs_101;
  wire [63:0] _result_T_103 = data_102 * coeffs_102;
  wire [63:0] _result_T_104 = data_103 * coeffs_103;
  wire [63:0] _result_T_105 = data_104 * coeffs_104;
  wire [63:0] _result_T_106 = data_105 * coeffs_105;
  wire [63:0] _result_T_107 = data_106 * coeffs_106;
  wire [63:0] _result_T_108 = data_107 * coeffs_107;
  wire [63:0] _result_T_109 = data_108 * coeffs_108;
  wire [63:0] _result_T_110 = data_109 * coeffs_109;
  wire [63:0] _result_T_111 = data_110 * coeffs_110;
  wire [63:0] _result_T_112 = data_111 * coeffs_111;
  wire [63:0] _result_T_113 = data_112 * coeffs_112;
  wire [63:0] _result_T_114 = data_113 * coeffs_113;
  wire [63:0] _result_T_115 = data_114 * coeffs_114;
  wire [63:0] _result_T_116 = data_115 * coeffs_115;
  wire [63:0] _result_T_117 = data_116 * coeffs_116;
  wire [63:0] _result_T_118 = data_117 * coeffs_117;
  wire [63:0] _result_T_119 = data_118 * coeffs_118;
  wire [63:0] _result_T_120 = data_119 * coeffs_119;
  wire [63:0] _result_T_121 = data_120 * coeffs_120;
  wire [63:0] _result_T_122 = data_121 * coeffs_121;
  wire [63:0] _result_T_123 = data_122 * coeffs_122;
  wire [63:0] _result_T_124 = data_123 * coeffs_123;
  wire [63:0] _result_T_125 = data_124 * coeffs_124;
  wire [63:0] _result_T_126 = data_125 * coeffs_125;
  wire [63:0] _result_T_127 = data_126 * coeffs_126;
  wire [63:0] _result_T_128 = data_127 * coeffs_127;
  wire [63:0] _result_T_129 = data_128 * coeffs_128;
  wire [63:0] _result_T_130 = data_129 * coeffs_129;
  wire [63:0] _result_T_131 = data_130 * coeffs_130;
  wire [63:0] _result_T_132 = data_131 * coeffs_131;
  wire [63:0] _result_T_133 = data_132 * coeffs_132;
  wire [63:0] _result_T_134 = data_133 * coeffs_133;
  wire [63:0] _result_T_135 = data_134 * coeffs_134;
  wire [63:0] _result_T_136 = data_135 * coeffs_135;
  wire [63:0] _result_T_137 = data_136 * coeffs_136;
  wire [63:0] _result_T_138 = data_137 * coeffs_137;
  wire [63:0] _result_T_139 = data_138 * coeffs_138;
  wire [63:0] _result_T_140 = data_139 * coeffs_139;
  wire [63:0] _result_T_141 = data_140 * coeffs_140;
  wire [63:0] _result_T_142 = data_141 * coeffs_141;
  wire [63:0] _result_T_143 = data_142 * coeffs_142;
  wire [63:0] _result_T_144 = data_143 * coeffs_143;
  wire [63:0] _result_T_145 = data_144 * coeffs_144;
  wire [63:0] _result_T_146 = data_145 * coeffs_145;
  wire [63:0] _result_T_147 = data_146 * coeffs_146;
  wire [63:0] _result_T_148 = data_147 * coeffs_147;
  wire [63:0] _result_T_149 = data_148 * coeffs_148;
  wire [63:0] _result_T_150 = data_149 * coeffs_149;
  wire [63:0] _result_T_151 = data_150 * coeffs_150;
  wire [63:0] _result_T_152 = data_151 * coeffs_151;
  wire [63:0] _result_T_153 = data_152 * coeffs_152;
  wire [63:0] _result_T_154 = data_153 * coeffs_153;
  wire [63:0] _result_T_155 = data_154 * coeffs_154;
  wire [63:0] _result_T_156 = data_155 * coeffs_155;
  wire [63:0] _result_T_157 = data_156 * coeffs_156;
  wire [63:0] _result_T_158 = data_157 * coeffs_157;
  wire [63:0] _result_T_159 = data_158 * coeffs_158;
  wire [63:0] _result_T_160 = data_159 * coeffs_159;
  wire [63:0] _result_T_161 = data_160 * coeffs_160;
  wire [63:0] _result_T_162 = data_161 * coeffs_161;
  wire [63:0] _result_T_163 = data_162 * coeffs_162;
  wire [63:0] _result_T_164 = data_163 * coeffs_163;
  wire [63:0] _result_T_165 = data_164 * coeffs_164;
  wire [63:0] _result_T_166 = data_165 * coeffs_165;
  wire [63:0] _result_T_167 = data_166 * coeffs_166;
  wire [63:0] _result_T_168 = data_167 * coeffs_167;
  wire [63:0] _result_T_169 = data_168 * coeffs_168;
  wire [63:0] _result_T_170 = data_169 * coeffs_169;
  wire [63:0] _result_T_171 = data_170 * coeffs_170;
  wire [63:0] _result_T_172 = data_171 * coeffs_171;
  wire [63:0] _result_T_173 = data_172 * coeffs_172;
  wire [63:0] _result_T_174 = data_173 * coeffs_173;
  wire [63:0] _result_T_175 = data_174 * coeffs_174;
  wire [63:0] _result_T_176 = data_175 * coeffs_175;
  wire [63:0] _result_T_177 = data_176 * coeffs_176;
  wire [63:0] _result_T_178 = data_177 * coeffs_177;
  wire [63:0] _result_T_179 = data_178 * coeffs_178;
  wire [63:0] _result_T_180 = data_179 * coeffs_179;
  wire [63:0] _result_T_181 = data_180 * coeffs_180;
  wire [63:0] _result_T_182 = data_181 * coeffs_181;
  wire [63:0] _result_T_183 = data_182 * coeffs_182;
  wire [63:0] _result_T_184 = data_183 * coeffs_183;
  wire [63:0] _result_T_185 = data_184 * coeffs_184;
  wire [63:0] _result_T_186 = data_185 * coeffs_185;
  wire [63:0] _result_T_187 = data_186 * coeffs_186;
  wire [63:0] _result_T_188 = data_187 * coeffs_187;
  wire [63:0] _result_T_189 = data_188 * coeffs_188;
  wire [63:0] _result_T_190 = data_189 * coeffs_189;
  wire [63:0] _result_T_191 = data_190 * coeffs_190;
  wire [63:0] _result_T_192 = data_191 * coeffs_191;
  wire [63:0] _result_T_193 = data_192 * coeffs_192;
  wire [63:0] _result_T_194 = data_193 * coeffs_193;
  wire [63:0] _result_T_195 = data_194 * coeffs_194;
  wire [63:0] _result_T_196 = data_195 * coeffs_195;
  wire [63:0] _result_T_197 = data_196 * coeffs_196;
  wire [63:0] _result_T_198 = data_197 * coeffs_197;
  wire [63:0] _result_T_199 = data_198 * coeffs_198;
  wire [63:0] _result_T_200 = data_199 * coeffs_199;
  wire [63:0] _result_T_201 = data_200 * coeffs_200;
  wire [63:0] _result_T_202 = data_201 * coeffs_201;
  wire [63:0] _result_T_203 = data_202 * coeffs_202;
  wire [63:0] _result_T_204 = data_203 * coeffs_203;
  wire [63:0] _result_T_205 = data_204 * coeffs_204;
  wire [63:0] _result_T_206 = data_205 * coeffs_205;
  wire [63:0] _result_T_207 = data_206 * coeffs_206;
  wire [63:0] _result_T_208 = data_207 * coeffs_207;
  wire [63:0] _result_T_209 = data_208 * coeffs_208;
  wire [63:0] _result_T_210 = data_209 * coeffs_209;
  wire [63:0] _result_T_211 = data_210 * coeffs_210;
  wire [63:0] _result_T_212 = data_211 * coeffs_211;
  wire [63:0] _result_T_213 = data_212 * coeffs_212;
  wire [63:0] _result_T_214 = data_213 * coeffs_213;
  wire [63:0] _result_T_215 = data_214 * coeffs_214;
  wire [63:0] _result_T_216 = data_215 * coeffs_215;
  wire [63:0] _result_T_217 = data_216 * coeffs_216;
  wire [63:0] _result_T_218 = data_217 * coeffs_217;
  wire [63:0] _result_T_219 = data_218 * coeffs_218;
  wire [63:0] _result_T_220 = data_219 * coeffs_219;
  wire [63:0] _result_T_221 = data_220 * coeffs_220;
  wire [63:0] _result_T_222 = data_221 * coeffs_221;
  wire [63:0] _result_T_223 = data_222 * coeffs_222;
  wire [63:0] _result_T_224 = data_223 * coeffs_223;
  wire [63:0] _result_T_225 = data_224 * coeffs_224;
  wire [63:0] _result_T_226 = data_225 * coeffs_225;
  wire [63:0] _result_T_227 = data_226 * coeffs_226;
  wire [63:0] _result_T_228 = data_227 * coeffs_227;
  wire [63:0] _result_T_229 = data_228 * coeffs_228;
  wire [63:0] _result_T_230 = data_229 * coeffs_229;
  wire [63:0] _result_T_231 = data_230 * coeffs_230;
  wire [63:0] _result_T_232 = data_231 * coeffs_231;
  wire [63:0] _result_T_233 = data_232 * coeffs_232;
  wire [63:0] _result_T_234 = data_233 * coeffs_233;
  wire [63:0] _result_T_235 = data_234 * coeffs_234;
  wire [63:0] _result_T_236 = data_235 * coeffs_235;
  wire [63:0] _result_T_237 = data_236 * coeffs_236;
  wire [63:0] _result_T_238 = data_237 * coeffs_237;
  wire [63:0] _result_T_239 = data_238 * coeffs_238;
  wire [63:0] _result_T_240 = data_239 * coeffs_239;
  wire [63:0] _result_T_241 = data_240 * coeffs_240;
  wire [63:0] _result_T_242 = data_241 * coeffs_241;
  wire [63:0] _result_T_243 = data_242 * coeffs_242;
  wire [63:0] _result_T_244 = data_243 * coeffs_243;
  wire [63:0] _result_T_245 = data_244 * coeffs_244;
  wire [63:0] _result_T_246 = data_245 * coeffs_245;
  wire [63:0] _result_T_247 = data_246 * coeffs_246;
  wire [63:0] _result_T_248 = data_247 * coeffs_247;
  wire [63:0] _result_T_249 = data_248 * coeffs_248;
  wire [63:0] _result_T_250 = data_249 * coeffs_249;
  wire [63:0] _result_T_251 = data_250 * coeffs_250;
  wire [63:0] _result_T_252 = data_251 * coeffs_251;
  wire [63:0] _result_T_253 = data_252 * coeffs_252;
  wire [63:0] _result_T_254 = data_253 * coeffs_253;
  wire [63:0] _result_T_255 = data_254 * coeffs_254;
  wire [63:0] _result_T_256 = data_255 * coeffs_255;
  wire [63:0] _result_T_257 = data_256 * coeffs_256;
  wire [63:0] _result_T_258 = data_257 * coeffs_257;
  wire [63:0] _result_T_259 = data_258 * coeffs_258;
  wire [63:0] _result_T_260 = data_259 * coeffs_259;
  wire [63:0] _result_T_261 = data_260 * coeffs_260;
  wire [63:0] _result_T_262 = data_261 * coeffs_261;
  wire [63:0] _result_T_263 = data_262 * coeffs_262;
  wire [63:0] _result_T_264 = data_263 * coeffs_263;
  wire [63:0] _result_T_265 = data_264 * coeffs_264;
  wire [63:0] _result_T_266 = data_265 * coeffs_265;
  wire [63:0] _result_T_267 = data_266 * coeffs_266;
  wire [63:0] _result_T_268 = data_267 * coeffs_267;
  wire [63:0] _result_T_269 = data_268 * coeffs_268;
  wire [63:0] _result_T_270 = data_269 * coeffs_269;
  wire [63:0] _result_T_271 = data_270 * coeffs_270;
  wire [63:0] _result_T_272 = data_271 * coeffs_271;
  wire [63:0] _result_T_273 = data_272 * coeffs_272;
  wire [63:0] _result_T_274 = data_273 * coeffs_273;
  wire [63:0] _result_T_275 = data_274 * coeffs_274;
  wire [63:0] _result_T_276 = data_275 * coeffs_275;
  wire [63:0] _result_T_277 = data_276 * coeffs_276;
  wire [63:0] _result_T_278 = data_277 * coeffs_277;
  wire [63:0] _result_T_279 = data_278 * coeffs_278;
  wire [63:0] _result_T_280 = data_279 * coeffs_279;
  wire [63:0] _result_T_281 = data_280 * coeffs_280;
  wire [63:0] _result_T_282 = data_281 * coeffs_281;
  wire [63:0] _result_T_283 = data_282 * coeffs_282;
  wire [63:0] _result_T_284 = data_283 * coeffs_283;
  wire [63:0] _result_T_285 = data_284 * coeffs_284;
  wire [63:0] _result_T_286 = data_285 * coeffs_285;
  wire [63:0] _result_T_287 = data_286 * coeffs_286;
  wire [63:0] _result_T_288 = data_287 * coeffs_287;
  wire [63:0] _result_T_289 = data_288 * coeffs_288;
  wire [63:0] _result_T_290 = data_289 * coeffs_289;
  wire [63:0] _result_T_291 = data_290 * coeffs_290;
  wire [63:0] _result_T_292 = data_291 * coeffs_291;
  wire [63:0] _result_T_293 = data_292 * coeffs_292;
  wire [63:0] _result_T_294 = data_293 * coeffs_293;
  wire [63:0] _result_T_295 = data_294 * coeffs_294;
  wire [63:0] _result_T_296 = data_295 * coeffs_295;
  wire [63:0] _result_T_297 = data_296 * coeffs_296;
  wire [63:0] _result_T_298 = data_297 * coeffs_297;
  wire [63:0] _result_T_299 = data_298 * coeffs_298;
  wire [63:0] _result_T_300 = data_299 * coeffs_299;
  wire [63:0] _result_T_301 = data_300 * coeffs_300;
  wire [63:0] _result_T_302 = data_301 * coeffs_301;
  wire [63:0] _result_T_303 = data_302 * coeffs_302;
  wire [63:0] _result_T_304 = data_303 * coeffs_303;
  wire [63:0] _result_T_305 = data_304 * coeffs_304;
  wire [63:0] _result_T_306 = data_305 * coeffs_305;
  wire [63:0] _result_T_307 = data_306 * coeffs_306;
  wire [63:0] _result_T_308 = data_307 * coeffs_307;
  wire [63:0] _result_T_309 = data_308 * coeffs_308;
  wire [63:0] _result_T_310 = data_309 * coeffs_309;
  wire [63:0] _result_T_311 = data_310 * coeffs_310;
  wire [63:0] _result_T_312 = data_311 * coeffs_311;
  wire [63:0] _result_T_313 = data_312 * coeffs_312;
  wire [63:0] _result_T_314 = data_313 * coeffs_313;
  wire [63:0] _result_T_315 = data_314 * coeffs_314;
  wire [63:0] _result_T_316 = data_315 * coeffs_315;
  wire [63:0] _result_T_317 = data_316 * coeffs_316;
  wire [63:0] _result_T_318 = data_317 * coeffs_317;
  wire [63:0] _result_T_319 = data_318 * coeffs_318;
  wire [63:0] _result_T_320 = data_319 * coeffs_319;
  wire [63:0] _result_T_321 = data_320 * coeffs_320;
  wire [63:0] _result_T_322 = data_321 * coeffs_321;
  wire [63:0] _result_T_323 = data_322 * coeffs_322;
  wire [63:0] _result_T_324 = data_323 * coeffs_323;
  wire [63:0] _result_T_325 = data_324 * coeffs_324;
  wire [63:0] _result_T_326 = data_325 * coeffs_325;
  wire [63:0] _result_T_327 = data_326 * coeffs_326;
  wire [63:0] _result_T_328 = data_327 * coeffs_327;
  wire [63:0] _result_T_329 = data_328 * coeffs_328;
  wire [63:0] _result_T_330 = data_329 * coeffs_329;
  wire [63:0] _result_T_331 = data_330 * coeffs_330;
  wire [63:0] _result_T_332 = data_331 * coeffs_331;
  wire [63:0] _result_T_333 = data_332 * coeffs_332;
  wire [63:0] _result_T_334 = data_333 * coeffs_333;
  wire [63:0] _result_T_335 = data_334 * coeffs_334;
  wire [63:0] _result_T_336 = data_335 * coeffs_335;
  wire [63:0] _result_T_337 = data_336 * coeffs_336;
  wire [63:0] _result_T_338 = data_337 * coeffs_337;
  wire [63:0] _result_T_339 = data_338 * coeffs_338;
  wire [63:0] _result_T_340 = data_339 * coeffs_339;
  wire [63:0] _result_T_341 = data_340 * coeffs_340;
  wire [63:0] _result_T_342 = data_341 * coeffs_341;
  wire [63:0] _result_T_343 = data_342 * coeffs_342;
  wire [63:0] _result_T_344 = data_343 * coeffs_343;
  wire [63:0] _result_T_345 = data_344 * coeffs_344;
  wire [63:0] _result_T_346 = data_345 * coeffs_345;
  wire [63:0] _result_T_347 = data_346 * coeffs_346;
  wire [63:0] _result_T_348 = data_347 * coeffs_347;
  wire [63:0] _result_T_349 = data_348 * coeffs_348;
  wire [63:0] _result_T_350 = data_349 * coeffs_349;
  wire [63:0] _result_T_351 = data_350 * coeffs_350;
  wire [63:0] _result_T_352 = data_351 * coeffs_351;
  wire [63:0] _result_T_353 = data_352 * coeffs_352;
  wire [63:0] _result_T_354 = data_353 * coeffs_353;
  wire [63:0] _result_T_355 = data_354 * coeffs_354;
  wire [63:0] _result_T_356 = data_355 * coeffs_355;
  wire [63:0] _result_T_357 = data_356 * coeffs_356;
  wire [63:0] _result_T_358 = data_357 * coeffs_357;
  wire [63:0] _result_T_359 = data_358 * coeffs_358;
  wire [63:0] _result_T_360 = data_359 * coeffs_359;
  wire [63:0] _result_T_361 = data_360 * coeffs_360;
  wire [63:0] _result_T_362 = data_361 * coeffs_361;
  wire [63:0] _result_T_363 = data_362 * coeffs_362;
  wire [63:0] _result_T_364 = data_363 * coeffs_363;
  wire [63:0] _result_T_365 = data_364 * coeffs_364;
  wire [63:0] _result_T_366 = data_365 * coeffs_365;
  wire [63:0] _result_T_367 = data_366 * coeffs_366;
  wire [63:0] _result_T_368 = data_367 * coeffs_367;
  wire [63:0] _result_T_369 = data_368 * coeffs_368;
  wire [63:0] _result_T_370 = data_369 * coeffs_369;
  wire [63:0] _result_T_371 = data_370 * coeffs_370;
  wire [63:0] _result_T_372 = data_371 * coeffs_371;
  wire [63:0] _result_T_373 = data_372 * coeffs_372;
  wire [63:0] _result_T_374 = data_373 * coeffs_373;
  wire [63:0] _result_T_375 = data_374 * coeffs_374;
  wire [63:0] _result_T_376 = data_375 * coeffs_375;
  wire [63:0] _result_T_377 = data_376 * coeffs_376;
  wire [63:0] _result_T_378 = data_377 * coeffs_377;
  wire [63:0] _result_T_379 = data_378 * coeffs_378;
  wire [63:0] _result_T_380 = data_379 * coeffs_379;
  wire [63:0] _result_T_381 = data_380 * coeffs_380;
  wire [63:0] _result_T_382 = data_381 * coeffs_381;
  wire [63:0] _result_T_383 = data_382 * coeffs_382;
  wire [63:0] _result_T_384 = data_383 * coeffs_383;
  wire [63:0] _result_T_385 = data_384 * coeffs_384;
  wire [63:0] _result_T_386 = data_385 * coeffs_385;
  wire [63:0] _result_T_387 = data_386 * coeffs_386;
  wire [63:0] _result_T_388 = data_387 * coeffs_387;
  wire [63:0] _result_T_389 = data_388 * coeffs_388;
  wire [63:0] _result_T_390 = data_389 * coeffs_389;
  wire [63:0] _result_T_391 = data_390 * coeffs_390;
  wire [63:0] _result_T_392 = data_391 * coeffs_391;
  wire [63:0] _result_T_393 = data_392 * coeffs_392;
  wire [63:0] _result_T_394 = data_393 * coeffs_393;
  wire [63:0] _result_T_395 = data_394 * coeffs_394;
  wire [63:0] _result_T_396 = data_395 * coeffs_395;
  wire [63:0] _result_T_397 = data_396 * coeffs_396;
  wire [63:0] _result_T_398 = data_397 * coeffs_397;
  wire [63:0] _result_T_399 = data_398 * coeffs_398;
  wire [63:0] _result_T_400 = data_399 * coeffs_399;
  wire [63:0] _result_T_401 = data_400 * coeffs_400;
  wire [63:0] _result_T_402 = data_401 * coeffs_401;
  wire [63:0] _result_T_403 = data_402 * coeffs_402;
  wire [63:0] _result_T_404 = data_403 * coeffs_403;
  wire [63:0] _result_T_405 = data_404 * coeffs_404;
  wire [63:0] _result_T_406 = data_405 * coeffs_405;
  wire [63:0] _result_T_407 = data_406 * coeffs_406;
  wire [63:0] _result_T_408 = data_407 * coeffs_407;
  wire [63:0] _result_T_409 = data_408 * coeffs_408;
  wire [63:0] _result_T_410 = data_409 * coeffs_409;
  wire [63:0] _result_T_411 = data_410 * coeffs_410;
  wire [63:0] _result_T_412 = data_411 * coeffs_411;
  wire [63:0] _result_T_413 = data_412 * coeffs_412;
  wire [63:0] _result_T_414 = data_413 * coeffs_413;
  wire [63:0] _result_T_415 = data_414 * coeffs_414;
  wire [63:0] _result_T_416 = data_415 * coeffs_415;
  wire [63:0] _result_T_417 = data_416 * coeffs_416;
  wire [63:0] _result_T_418 = data_417 * coeffs_417;
  wire [63:0] _result_T_419 = data_418 * coeffs_418;
  wire [63:0] _result_T_420 = data_419 * coeffs_419;
  wire [63:0] _result_T_421 = data_420 * coeffs_420;
  wire [63:0] _result_T_422 = data_421 * coeffs_421;
  wire [63:0] _result_T_423 = data_422 * coeffs_422;
  wire [63:0] _result_T_424 = data_423 * coeffs_423;
  wire [63:0] _result_T_425 = data_424 * coeffs_424;
  wire [63:0] _result_T_426 = data_425 * coeffs_425;
  wire [63:0] _result_T_427 = data_426 * coeffs_426;
  wire [63:0] _result_T_428 = data_427 * coeffs_427;
  wire [63:0] _result_T_429 = data_428 * coeffs_428;
  wire [63:0] _result_T_430 = data_429 * coeffs_429;
  wire [63:0] _result_T_431 = data_430 * coeffs_430;
  wire [63:0] _result_T_432 = data_431 * coeffs_431;
  wire [63:0] _result_T_433 = data_432 * coeffs_432;
  wire [63:0] _result_T_434 = data_433 * coeffs_433;
  wire [63:0] _result_T_435 = data_434 * coeffs_434;
  wire [63:0] _result_T_436 = data_435 * coeffs_435;
  wire [63:0] _result_T_437 = data_436 * coeffs_436;
  wire [63:0] _result_T_438 = data_437 * coeffs_437;
  wire [63:0] _result_T_439 = data_438 * coeffs_438;
  wire [63:0] _result_T_440 = data_439 * coeffs_439;
  wire [63:0] _result_T_441 = data_440 * coeffs_440;
  wire [63:0] _result_T_442 = data_441 * coeffs_441;
  wire [63:0] _result_T_443 = data_442 * coeffs_442;
  wire [63:0] _result_T_444 = data_443 * coeffs_443;
  wire [63:0] _result_T_445 = data_444 * coeffs_444;
  wire [63:0] _result_T_446 = data_445 * coeffs_445;
  wire [63:0] _result_T_447 = data_446 * coeffs_446;
  wire [63:0] _result_T_448 = data_447 * coeffs_447;
  wire [63:0] _result_T_449 = data_448 * coeffs_448;
  wire [63:0] _result_T_450 = data_449 * coeffs_449;
  wire [63:0] _result_T_451 = data_450 * coeffs_450;
  wire [63:0] _result_T_452 = data_451 * coeffs_451;
  wire [63:0] _result_T_453 = data_452 * coeffs_452;
  wire [63:0] _result_T_454 = data_453 * coeffs_453;
  wire [63:0] _result_T_455 = data_454 * coeffs_454;
  wire [63:0] _result_T_456 = data_455 * coeffs_455;
  wire [63:0] _result_T_457 = data_456 * coeffs_456;
  wire [63:0] _result_T_458 = data_457 * coeffs_457;
  wire [63:0] _result_T_459 = data_458 * coeffs_458;
  wire [63:0] _result_T_460 = data_459 * coeffs_459;
  wire [63:0] _result_T_461 = data_460 * coeffs_460;
  wire [63:0] _result_T_462 = data_461 * coeffs_461;
  wire [63:0] _result_T_463 = data_462 * coeffs_462;
  wire [63:0] _result_T_464 = data_463 * coeffs_463;
  wire [63:0] _result_T_465 = data_464 * coeffs_464;
  wire [63:0] _result_T_466 = data_465 * coeffs_465;
  wire [63:0] _result_T_467 = data_466 * coeffs_466;
  wire [63:0] _result_T_468 = data_467 * coeffs_467;
  wire [63:0] _result_T_469 = data_468 * coeffs_468;
  wire [63:0] _result_T_470 = data_469 * coeffs_469;
  wire [63:0] _result_T_471 = data_470 * coeffs_470;
  wire [63:0] _result_T_472 = data_471 * coeffs_471;
  wire [63:0] _result_T_473 = data_472 * coeffs_472;
  wire [63:0] _result_T_474 = data_473 * coeffs_473;
  wire [63:0] _result_T_475 = data_474 * coeffs_474;
  wire [63:0] _result_T_476 = data_475 * coeffs_475;
  wire [63:0] _result_T_477 = data_476 * coeffs_476;
  wire [63:0] _result_T_478 = data_477 * coeffs_477;
  wire [63:0] _result_T_479 = data_478 * coeffs_478;
  wire [63:0] _result_T_480 = data_479 * coeffs_479;
  wire [63:0] _result_T_481 = data_480 * coeffs_480;
  wire [63:0] _result_T_482 = data_481 * coeffs_481;
  wire [63:0] _result_T_483 = data_482 * coeffs_482;
  wire [63:0] _result_T_484 = data_483 * coeffs_483;
  wire [63:0] _result_T_485 = data_484 * coeffs_484;
  wire [63:0] _result_T_486 = data_485 * coeffs_485;
  wire [63:0] _result_T_487 = data_486 * coeffs_486;
  wire [63:0] _result_T_488 = data_487 * coeffs_487;
  wire [63:0] _result_T_489 = data_488 * coeffs_488;
  wire [63:0] _result_T_490 = data_489 * coeffs_489;
  wire [63:0] _result_T_491 = data_490 * coeffs_490;
  wire [63:0] _result_T_492 = data_491 * coeffs_491;
  wire [63:0] _result_T_493 = data_492 * coeffs_492;
  wire [63:0] _result_T_494 = data_493 * coeffs_493;
  wire [63:0] _result_T_495 = data_494 * coeffs_494;
  wire [63:0] _result_T_496 = data_495 * coeffs_495;
  wire [63:0] _result_T_497 = data_496 * coeffs_496;
  wire [63:0] _result_T_498 = data_497 * coeffs_497;
  wire [63:0] _result_T_499 = data_498 * coeffs_498;
  wire [63:0] _result_T_500 = data_499 * coeffs_499;
  wire [63:0] _result_T_501 = data_500 * coeffs_500;
  wire [63:0] _result_T_502 = data_501 * coeffs_501;
  wire [63:0] _result_T_503 = data_502 * coeffs_502;
  wire [63:0] _result_T_504 = data_503 * coeffs_503;
  wire [63:0] _result_T_505 = data_504 * coeffs_504;
  wire [63:0] _result_T_506 = data_505 * coeffs_505;
  wire [63:0] _result_T_507 = data_506 * coeffs_506;
  wire [63:0] _result_T_508 = data_507 * coeffs_507;
  wire [63:0] _result_T_509 = data_508 * coeffs_508;
  wire [63:0] _result_T_510 = data_509 * coeffs_509;
  wire [63:0] _result_T_511 = data_510 * coeffs_510;
  wire [63:0] _result_T_512 = data_511 * coeffs_511;
  wire [63:0] _result_T_513 = data_512 * coeffs_512;
  wire [63:0] _result_T_514 = data_513 * coeffs_513;
  wire [63:0] _result_T_515 = data_514 * coeffs_514;
  wire [63:0] _result_T_516 = data_515 * coeffs_515;
  wire [63:0] _result_T_517 = data_516 * coeffs_516;
  wire [63:0] _result_T_518 = data_517 * coeffs_517;
  wire [63:0] _result_T_519 = data_518 * coeffs_518;
  wire [63:0] _result_T_520 = data_519 * coeffs_519;
  wire [63:0] _result_T_521 = data_520 * coeffs_520;
  wire [63:0] _result_T_522 = data_521 * coeffs_521;
  wire [63:0] _result_T_523 = data_522 * coeffs_522;
  wire [63:0] _result_T_524 = data_523 * coeffs_523;
  wire [63:0] _result_T_525 = data_524 * coeffs_524;
  wire [63:0] _result_T_526 = data_525 * coeffs_525;
  wire [63:0] _result_T_527 = data_526 * coeffs_526;
  wire [63:0] _result_T_528 = data_527 * coeffs_527;
  wire [63:0] _result_T_529 = data_528 * coeffs_528;
  wire [63:0] _result_T_530 = data_529 * coeffs_529;
  wire [63:0] _result_T_531 = data_530 * coeffs_530;
  wire [63:0] _result_T_532 = data_531 * coeffs_531;
  wire [63:0] _result_T_533 = data_532 * coeffs_532;
  wire [63:0] _result_T_534 = data_533 * coeffs_533;
  wire [63:0] _result_T_535 = data_534 * coeffs_534;
  wire [63:0] _result_T_536 = data_535 * coeffs_535;
  wire [63:0] _result_T_537 = data_536 * coeffs_536;
  wire [63:0] _result_T_538 = data_537 * coeffs_537;
  wire [63:0] _result_T_539 = data_538 * coeffs_538;
  wire [63:0] _result_T_540 = data_539 * coeffs_539;
  wire [63:0] _result_T_541 = data_540 * coeffs_540;
  wire [63:0] _result_T_542 = data_541 * coeffs_541;
  wire [63:0] _result_T_543 = data_542 * coeffs_542;
  wire [63:0] _result_T_544 = data_543 * coeffs_543;
  wire [63:0] _result_T_545 = data_544 * coeffs_544;
  wire [63:0] _result_T_546 = data_545 * coeffs_545;
  wire [63:0] _result_T_547 = data_546 * coeffs_546;
  wire [63:0] _result_T_548 = data_547 * coeffs_547;
  wire [63:0] _result_T_549 = data_548 * coeffs_548;
  wire [63:0] _result_T_550 = data_549 * coeffs_549;
  wire [63:0] _result_T_551 = data_550 * coeffs_550;
  wire [63:0] _result_T_552 = data_551 * coeffs_551;
  wire [63:0] _result_T_553 = data_552 * coeffs_552;
  wire [63:0] _result_T_554 = data_553 * coeffs_553;
  wire [63:0] _result_T_555 = data_554 * coeffs_554;
  wire [63:0] _result_T_556 = data_555 * coeffs_555;
  wire [63:0] _result_T_557 = data_556 * coeffs_556;
  wire [63:0] _result_T_558 = data_557 * coeffs_557;
  wire [63:0] _result_T_559 = data_558 * coeffs_558;
  wire [63:0] _result_T_560 = data_559 * coeffs_559;
  wire [63:0] _result_T_561 = data_560 * coeffs_560;
  wire [63:0] _result_T_562 = data_561 * coeffs_561;
  wire [63:0] _result_T_563 = data_562 * coeffs_562;
  wire [63:0] _result_T_564 = data_563 * coeffs_563;
  wire [63:0] _result_T_565 = data_564 * coeffs_564;
  wire [63:0] _result_T_566 = data_565 * coeffs_565;
  wire [63:0] _result_T_567 = data_566 * coeffs_566;
  wire [63:0] _result_T_568 = data_567 * coeffs_567;
  wire [63:0] _result_T_569 = data_568 * coeffs_568;
  wire [63:0] _result_T_570 = data_569 * coeffs_569;
  wire [63:0] _result_T_571 = data_570 * coeffs_570;
  wire [63:0] _result_T_572 = data_571 * coeffs_571;
  wire [63:0] _result_T_573 = data_572 * coeffs_572;
  wire [63:0] _result_T_574 = data_573 * coeffs_573;
  wire [63:0] _result_T_575 = data_574 * coeffs_574;
  wire [63:0] _result_T_576 = data_575 * coeffs_575;
  wire [63:0] _result_T_577 = data_576 * coeffs_576;
  wire [63:0] _result_T_578 = data_577 * coeffs_577;
  wire [63:0] _result_T_579 = data_578 * coeffs_578;
  wire [63:0] _result_T_580 = data_579 * coeffs_579;
  wire [63:0] _result_T_581 = data_580 * coeffs_580;
  wire [63:0] _result_T_582 = data_581 * coeffs_581;
  wire [63:0] _result_T_583 = data_582 * coeffs_582;
  wire [63:0] _result_T_584 = data_583 * coeffs_583;
  wire [63:0] _result_T_585 = data_584 * coeffs_584;
  wire [63:0] _result_T_586 = data_585 * coeffs_585;
  wire [63:0] _result_T_587 = data_586 * coeffs_586;
  wire [63:0] _result_T_588 = data_587 * coeffs_587;
  wire [63:0] _result_T_589 = data_588 * coeffs_588;
  wire [63:0] _result_T_590 = data_589 * coeffs_589;
  wire [63:0] _result_T_591 = data_590 * coeffs_590;
  wire [63:0] _result_T_592 = data_591 * coeffs_591;
  wire [63:0] _result_T_593 = data_592 * coeffs_592;
  wire [63:0] _result_T_594 = data_593 * coeffs_593;
  wire [63:0] _result_T_595 = data_594 * coeffs_594;
  wire [63:0] _result_T_596 = data_595 * coeffs_595;
  wire [63:0] _result_T_597 = data_596 * coeffs_596;
  wire [63:0] _result_T_598 = data_597 * coeffs_597;
  wire [63:0] _result_T_599 = data_598 * coeffs_598;
  wire [63:0] _result_T_600 = data_599 * coeffs_599;
  wire [63:0] _result_T_601 = data_600 * coeffs_600;
  wire [63:0] _result_T_602 = data_601 * coeffs_601;
  wire [63:0] _result_T_603 = data_602 * coeffs_602;
  wire [63:0] _result_T_604 = data_603 * coeffs_603;
  wire [63:0] _result_T_605 = data_604 * coeffs_604;
  wire [63:0] _result_T_606 = data_605 * coeffs_605;
  wire [63:0] _result_T_607 = data_606 * coeffs_606;
  wire [63:0] _result_T_608 = data_607 * coeffs_607;
  wire [63:0] _result_T_609 = data_608 * coeffs_608;
  wire [63:0] _result_T_610 = data_609 * coeffs_609;
  wire [63:0] _result_T_611 = data_610 * coeffs_610;
  wire [63:0] _result_T_612 = data_611 * coeffs_611;
  wire [63:0] _result_T_613 = data_612 * coeffs_612;
  wire [63:0] _result_T_614 = data_613 * coeffs_613;
  wire [63:0] _result_T_615 = data_614 * coeffs_614;
  wire [63:0] _result_T_616 = data_615 * coeffs_615;
  wire [63:0] _result_T_617 = data_616 * coeffs_616;
  wire [63:0] _result_T_618 = data_617 * coeffs_617;
  wire [63:0] _result_T_619 = data_618 * coeffs_618;
  wire [63:0] _result_T_620 = data_619 * coeffs_619;
  wire [63:0] _result_T_621 = data_620 * coeffs_620;
  wire [63:0] _result_T_622 = data_621 * coeffs_621;
  wire [63:0] _result_T_623 = data_622 * coeffs_622;
  wire [63:0] _result_T_624 = data_623 * coeffs_623;
  wire [63:0] _result_T_625 = data_624 * coeffs_624;
  wire [63:0] _result_T_626 = data_625 * coeffs_625;
  wire [63:0] _result_T_627 = data_626 * coeffs_626;
  wire [63:0] _result_T_628 = data_627 * coeffs_627;
  wire [63:0] _result_T_629 = data_628 * coeffs_628;
  wire [63:0] _result_T_630 = data_629 * coeffs_629;
  wire [63:0] _result_T_631 = data_630 * coeffs_630;
  wire [63:0] _result_T_632 = data_631 * coeffs_631;
  wire [63:0] _result_T_633 = data_632 * coeffs_632;
  wire [63:0] _result_T_634 = data_633 * coeffs_633;
  wire [63:0] _result_T_635 = data_634 * coeffs_634;
  wire [63:0] _result_T_636 = data_635 * coeffs_635;
  wire [63:0] _result_T_637 = data_636 * coeffs_636;
  wire [63:0] _result_T_638 = data_637 * coeffs_637;
  wire [63:0] _result_T_639 = data_638 * coeffs_638;
  wire [63:0] _result_T_640 = data_639 * coeffs_639;
  wire [63:0] _result_T_641 = data_640 * coeffs_640;
  wire [63:0] _result_T_642 = data_641 * coeffs_641;
  wire [63:0] _result_T_643 = data_642 * coeffs_642;
  wire [63:0] _result_T_644 = data_643 * coeffs_643;
  wire [63:0] _result_T_645 = data_644 * coeffs_644;
  wire [63:0] _result_T_646 = data_645 * coeffs_645;
  wire [63:0] _result_T_647 = data_646 * coeffs_646;
  wire [63:0] _result_T_648 = data_647 * coeffs_647;
  wire [63:0] _result_T_649 = data_648 * coeffs_648;
  wire [63:0] _result_T_650 = data_649 * coeffs_649;
  wire [63:0] _result_T_651 = data_650 * coeffs_650;
  wire [63:0] _result_T_652 = data_651 * coeffs_651;
  wire [63:0] _result_T_653 = data_652 * coeffs_652;
  wire [63:0] _result_T_654 = data_653 * coeffs_653;
  wire [63:0] _result_T_655 = data_654 * coeffs_654;
  wire [63:0] _result_T_656 = data_655 * coeffs_655;
  wire [63:0] _result_T_657 = data_656 * coeffs_656;
  wire [63:0] _result_T_658 = data_657 * coeffs_657;
  wire [63:0] _result_T_659 = data_658 * coeffs_658;
  wire [63:0] _result_T_660 = data_659 * coeffs_659;
  wire [63:0] _result_T_661 = data_660 * coeffs_660;
  wire [63:0] _result_T_662 = data_661 * coeffs_661;
  wire [63:0] _result_T_663 = data_662 * coeffs_662;
  wire [63:0] _result_T_664 = data_663 * coeffs_663;
  wire [63:0] _result_T_665 = data_664 * coeffs_664;
  wire [63:0] _result_T_666 = data_665 * coeffs_665;
  wire [63:0] _result_T_667 = data_666 * coeffs_666;
  wire [63:0] _result_T_668 = data_667 * coeffs_667;
  wire [63:0] _result_T_669 = data_668 * coeffs_668;
  wire [63:0] _result_T_670 = data_669 * coeffs_669;
  wire [63:0] _result_T_671 = data_670 * coeffs_670;
  wire [63:0] _result_T_672 = data_671 * coeffs_671;
  wire [63:0] _result_T_673 = data_672 * coeffs_672;
  wire [63:0] _result_T_674 = data_673 * coeffs_673;
  wire [63:0] _result_T_675 = data_674 * coeffs_674;
  wire [63:0] _result_T_676 = data_675 * coeffs_675;
  wire [63:0] _result_T_677 = data_676 * coeffs_676;
  wire [63:0] _result_T_678 = data_677 * coeffs_677;
  wire [63:0] _result_T_679 = data_678 * coeffs_678;
  wire [63:0] _result_T_680 = data_679 * coeffs_679;
  wire [63:0] _result_T_681 = data_680 * coeffs_680;
  wire [63:0] _result_T_682 = data_681 * coeffs_681;
  wire [63:0] _result_T_683 = data_682 * coeffs_682;
  wire [63:0] _result_T_684 = data_683 * coeffs_683;
  wire [63:0] _result_T_685 = data_684 * coeffs_684;
  wire [63:0] _result_T_686 = data_685 * coeffs_685;
  wire [63:0] _result_T_687 = data_686 * coeffs_686;
  wire [63:0] _result_T_688 = data_687 * coeffs_687;
  wire [63:0] _result_T_689 = data_688 * coeffs_688;
  wire [63:0] _result_T_690 = data_689 * coeffs_689;
  wire [63:0] _result_T_691 = data_690 * coeffs_690;
  wire [63:0] _result_T_692 = data_691 * coeffs_691;
  wire [63:0] _result_T_693 = data_692 * coeffs_692;
  wire [63:0] _result_T_694 = data_693 * coeffs_693;
  wire [63:0] _result_T_695 = data_694 * coeffs_694;
  wire [63:0] _result_T_696 = data_695 * coeffs_695;
  wire [63:0] _result_T_697 = data_696 * coeffs_696;
  wire [63:0] _result_T_698 = data_697 * coeffs_697;
  wire [63:0] _result_T_699 = data_698 * coeffs_698;
  wire [63:0] _result_T_700 = data_699 * coeffs_699;
  wire [63:0] _result_T_701 = data_700 * coeffs_700;
  wire [63:0] _result_T_702 = data_701 * coeffs_701;
  wire [63:0] _result_T_703 = data_702 * coeffs_702;
  wire [63:0] _result_T_704 = data_703 * coeffs_703;
  wire [63:0] _result_T_705 = data_704 * coeffs_704;
  wire [63:0] _result_T_706 = data_705 * coeffs_705;
  wire [63:0] _result_T_707 = data_706 * coeffs_706;
  wire [63:0] _result_T_708 = data_707 * coeffs_707;
  wire [63:0] _result_T_709 = data_708 * coeffs_708;
  wire [63:0] _result_T_710 = data_709 * coeffs_709;
  wire [63:0] _result_T_711 = data_710 * coeffs_710;
  wire [63:0] _result_T_712 = data_711 * coeffs_711;
  wire [63:0] _result_T_713 = data_712 * coeffs_712;
  wire [63:0] _result_T_714 = data_713 * coeffs_713;
  wire [63:0] _result_T_715 = data_714 * coeffs_714;
  wire [63:0] _result_T_716 = data_715 * coeffs_715;
  wire [63:0] _result_T_717 = data_716 * coeffs_716;
  wire [63:0] _result_T_718 = data_717 * coeffs_717;
  wire [63:0] _result_T_719 = data_718 * coeffs_718;
  wire [63:0] _result_T_720 = data_719 * coeffs_719;
  wire [63:0] _result_T_721 = data_720 * coeffs_720;
  wire [63:0] _result_T_722 = data_721 * coeffs_721;
  wire [63:0] _result_T_723 = data_722 * coeffs_722;
  wire [63:0] _result_T_724 = data_723 * coeffs_723;
  wire [63:0] _result_T_725 = data_724 * coeffs_724;
  wire [63:0] _result_T_726 = data_725 * coeffs_725;
  wire [63:0] _result_T_727 = data_726 * coeffs_726;
  wire [63:0] _result_T_728 = data_727 * coeffs_727;
  wire [63:0] _result_T_729 = data_728 * coeffs_728;
  wire [63:0] _result_T_730 = data_729 * coeffs_729;
  wire [63:0] _result_T_731 = data_730 * coeffs_730;
  wire [63:0] _result_T_732 = data_731 * coeffs_731;
  wire [63:0] _result_T_733 = data_732 * coeffs_732;
  wire [63:0] _result_T_734 = data_733 * coeffs_733;
  wire [63:0] _result_T_735 = data_734 * coeffs_734;
  wire [63:0] _result_T_736 = data_735 * coeffs_735;
  wire [63:0] _result_T_737 = data_736 * coeffs_736;
  wire [63:0] _result_T_738 = data_737 * coeffs_737;
  wire [63:0] _result_T_739 = data_738 * coeffs_738;
  wire [63:0] _result_T_740 = data_739 * coeffs_739;
  wire [63:0] _result_T_741 = data_740 * coeffs_740;
  wire [63:0] _result_T_742 = data_741 * coeffs_741;
  wire [63:0] _result_T_743 = data_742 * coeffs_742;
  wire [63:0] _result_T_744 = data_743 * coeffs_743;
  wire [63:0] _result_T_745 = data_744 * coeffs_744;
  wire [63:0] _result_T_746 = data_745 * coeffs_745;
  wire [63:0] _result_T_747 = data_746 * coeffs_746;
  wire [63:0] _result_T_748 = data_747 * coeffs_747;
  wire [63:0] _result_T_749 = data_748 * coeffs_748;
  wire [63:0] _result_T_750 = data_749 * coeffs_749;
  wire [63:0] _result_T_751 = data_750 * coeffs_750;
  wire [63:0] _result_T_752 = data_751 * coeffs_751;
  wire [63:0] _result_T_753 = data_752 * coeffs_752;
  wire [63:0] _result_T_754 = data_753 * coeffs_753;
  wire [63:0] _result_T_755 = data_754 * coeffs_754;
  wire [63:0] _result_T_756 = data_755 * coeffs_755;
  wire [63:0] _result_T_757 = data_756 * coeffs_756;
  wire [63:0] _result_T_758 = data_757 * coeffs_757;
  wire [63:0] _result_T_759 = data_758 * coeffs_758;
  wire [63:0] _result_T_760 = data_759 * coeffs_759;
  wire [63:0] _result_T_761 = data_760 * coeffs_760;
  wire [63:0] _result_T_762 = data_761 * coeffs_761;
  wire [63:0] _result_T_763 = data_762 * coeffs_762;
  wire [63:0] _result_T_764 = data_763 * coeffs_763;
  wire [63:0] _result_T_765 = data_764 * coeffs_764;
  wire [63:0] _result_T_766 = data_765 * coeffs_765;
  wire [63:0] _result_T_767 = data_766 * coeffs_766;
  wire [63:0] _result_T_768 = data_767 * coeffs_767;
  wire [63:0] _result_T_769 = data_768 * coeffs_768;
  wire [63:0] _result_T_770 = data_769 * coeffs_769;
  wire [63:0] _result_T_771 = data_770 * coeffs_770;
  wire [63:0] _result_T_772 = data_771 * coeffs_771;
  wire [63:0] _result_T_773 = data_772 * coeffs_772;
  wire [63:0] _result_T_774 = data_773 * coeffs_773;
  wire [63:0] _result_T_775 = data_774 * coeffs_774;
  wire [63:0] _result_T_776 = data_775 * coeffs_775;
  wire [63:0] _result_T_777 = data_776 * coeffs_776;
  wire [63:0] _result_T_778 = data_777 * coeffs_777;
  wire [63:0] _result_T_779 = data_778 * coeffs_778;
  wire [63:0] _result_T_780 = data_779 * coeffs_779;
  wire [63:0] _result_T_781 = data_780 * coeffs_780;
  wire [63:0] _result_T_782 = data_781 * coeffs_781;
  wire [63:0] _result_T_783 = data_782 * coeffs_782;
  wire [63:0] _result_T_784 = data_783 * coeffs_783;
  wire [63:0] _result_T_785 = data_784 * coeffs_784;
  wire [63:0] _result_T_786 = data_785 * coeffs_785;
  wire [63:0] _result_T_787 = data_786 * coeffs_786;
  wire [63:0] _result_T_788 = data_787 * coeffs_787;
  wire [63:0] _result_T_789 = data_788 * coeffs_788;
  wire [63:0] _result_T_790 = data_789 * coeffs_789;
  wire [63:0] _result_T_791 = data_790 * coeffs_790;
  wire [63:0] _result_T_792 = data_791 * coeffs_791;
  wire [63:0] _result_T_793 = data_792 * coeffs_792;
  wire [63:0] _result_T_794 = data_793 * coeffs_793;
  wire [63:0] _result_T_795 = data_794 * coeffs_794;
  wire [63:0] _result_T_796 = data_795 * coeffs_795;
  wire [63:0] _result_T_797 = data_796 * coeffs_796;
  wire [63:0] _result_T_798 = data_797 * coeffs_797;
  wire [63:0] _result_T_799 = data_798 * coeffs_798;
  wire [63:0] _result_T_800 = data_799 * coeffs_799;
  wire [63:0] _result_T_801 = data_800 * coeffs_800;
  wire [63:0] _result_T_802 = data_801 * coeffs_801;
  wire [63:0] _result_T_803 = data_802 * coeffs_802;
  wire [63:0] _result_T_804 = data_803 * coeffs_803;
  wire [63:0] _result_T_805 = data_804 * coeffs_804;
  wire [63:0] _result_T_806 = data_805 * coeffs_805;
  wire [63:0] _result_T_807 = data_806 * coeffs_806;
  wire [63:0] _result_T_808 = data_807 * coeffs_807;
  wire [63:0] _result_T_809 = data_808 * coeffs_808;
  wire [63:0] _result_T_810 = data_809 * coeffs_809;
  wire [63:0] _result_T_811 = data_810 * coeffs_810;
  wire [63:0] _result_T_812 = data_811 * coeffs_811;
  wire [63:0] _result_T_813 = data_812 * coeffs_812;
  wire [63:0] _result_T_814 = data_813 * coeffs_813;
  wire [63:0] _result_T_815 = data_814 * coeffs_814;
  wire [63:0] _result_T_816 = data_815 * coeffs_815;
  wire [63:0] _result_T_817 = data_816 * coeffs_816;
  wire [63:0] _result_T_818 = data_817 * coeffs_817;
  wire [63:0] _result_T_819 = data_818 * coeffs_818;
  wire [63:0] _result_T_820 = data_819 * coeffs_819;
  wire [63:0] _result_T_821 = data_820 * coeffs_820;
  wire [63:0] _result_T_822 = data_821 * coeffs_821;
  wire [63:0] _result_T_823 = data_822 * coeffs_822;
  wire [63:0] _result_T_824 = data_823 * coeffs_823;
  wire [63:0] _result_T_825 = data_824 * coeffs_824;
  wire [63:0] _result_T_826 = data_825 * coeffs_825;
  wire [63:0] _result_T_827 = data_826 * coeffs_826;
  wire [63:0] _result_T_828 = data_827 * coeffs_827;
  wire [63:0] _result_T_829 = data_828 * coeffs_828;
  wire [63:0] _result_T_830 = data_829 * coeffs_829;
  wire [63:0] _result_T_831 = data_830 * coeffs_830;
  wire [63:0] _result_T_832 = data_831 * coeffs_831;
  wire [63:0] _result_T_833 = data_832 * coeffs_832;
  wire [63:0] _result_T_834 = data_833 * coeffs_833;
  wire [63:0] _result_T_835 = data_834 * coeffs_834;
  wire [63:0] _result_T_836 = data_835 * coeffs_835;
  wire [63:0] _result_T_837 = data_836 * coeffs_836;
  wire [63:0] _result_T_838 = data_837 * coeffs_837;
  wire [63:0] _result_T_839 = data_838 * coeffs_838;
  wire [63:0] _result_T_840 = data_839 * coeffs_839;
  wire [63:0] _result_T_841 = data_840 * coeffs_840;
  wire [63:0] _result_T_842 = data_841 * coeffs_841;
  wire [63:0] _result_T_843 = data_842 * coeffs_842;
  wire [63:0] _result_T_844 = data_843 * coeffs_843;
  wire [63:0] _result_T_845 = data_844 * coeffs_844;
  wire [63:0] _result_T_846 = data_845 * coeffs_845;
  wire [63:0] _result_T_847 = data_846 * coeffs_846;
  wire [63:0] _result_T_848 = data_847 * coeffs_847;
  wire [63:0] _result_T_849 = data_848 * coeffs_848;
  wire [63:0] _result_T_850 = data_849 * coeffs_849;
  wire [63:0] _result_T_851 = data_850 * coeffs_850;
  wire [63:0] _result_T_852 = data_851 * coeffs_851;
  wire [63:0] _result_T_853 = data_852 * coeffs_852;
  wire [63:0] _result_T_854 = data_853 * coeffs_853;
  wire [63:0] _result_T_855 = data_854 * coeffs_854;
  wire [63:0] _result_T_856 = data_855 * coeffs_855;
  wire [63:0] _result_T_857 = data_856 * coeffs_856;
  wire [63:0] _result_T_858 = data_857 * coeffs_857;
  wire [63:0] _result_T_859 = data_858 * coeffs_858;
  wire [63:0] _result_T_860 = data_859 * coeffs_859;
  wire [63:0] _result_T_861 = data_860 * coeffs_860;
  wire [63:0] _result_T_862 = data_861 * coeffs_861;
  wire [63:0] _result_T_863 = data_862 * coeffs_862;
  wire [63:0] _result_T_864 = data_863 * coeffs_863;
  wire [63:0] _result_T_865 = data_864 * coeffs_864;
  wire [63:0] _result_T_866 = data_865 * coeffs_865;
  wire [63:0] _result_T_867 = data_866 * coeffs_866;
  wire [63:0] _result_T_868 = data_867 * coeffs_867;
  wire [63:0] _result_T_869 = data_868 * coeffs_868;
  wire [63:0] _result_T_870 = data_869 * coeffs_869;
  wire [63:0] _result_T_871 = data_870 * coeffs_870;
  wire [63:0] _result_T_872 = data_871 * coeffs_871;
  wire [63:0] _result_T_873 = data_872 * coeffs_872;
  wire [63:0] _result_T_874 = data_873 * coeffs_873;
  wire [63:0] _result_T_875 = data_874 * coeffs_874;
  wire [63:0] _result_T_876 = data_875 * coeffs_875;
  wire [63:0] _result_T_877 = data_876 * coeffs_876;
  wire [63:0] _result_T_878 = data_877 * coeffs_877;
  wire [63:0] _result_T_879 = data_878 * coeffs_878;
  wire [63:0] _result_T_880 = data_879 * coeffs_879;
  wire [63:0] _result_T_881 = data_880 * coeffs_880;
  wire [63:0] _result_T_882 = data_881 * coeffs_881;
  wire [63:0] _result_T_883 = data_882 * coeffs_882;
  wire [63:0] _result_T_884 = data_883 * coeffs_883;
  wire [63:0] _result_T_885 = data_884 * coeffs_884;
  wire [63:0] _result_T_886 = data_885 * coeffs_885;
  wire [63:0] _result_T_887 = data_886 * coeffs_886;
  wire [63:0] _result_T_888 = data_887 * coeffs_887;
  wire [63:0] _result_T_889 = data_888 * coeffs_888;
  wire [63:0] _result_T_890 = data_889 * coeffs_889;
  wire [63:0] _result_T_891 = data_890 * coeffs_890;
  wire [63:0] _result_T_892 = data_891 * coeffs_891;
  wire [63:0] _result_T_893 = data_892 * coeffs_892;
  wire [63:0] _result_T_894 = data_893 * coeffs_893;
  wire [63:0] _result_T_895 = data_894 * coeffs_894;
  wire [63:0] _result_T_896 = data_895 * coeffs_895;
  wire [63:0] _result_T_897 = data_896 * coeffs_896;
  wire [63:0] _result_T_898 = data_897 * coeffs_897;
  wire [63:0] _result_T_899 = data_898 * coeffs_898;
  wire [63:0] _result_T_900 = data_899 * coeffs_899;
  wire [63:0] _result_T_901 = data_900 * coeffs_900;
  wire [63:0] _result_T_902 = data_901 * coeffs_901;
  wire [63:0] _result_T_903 = data_902 * coeffs_902;
  wire [63:0] _result_T_904 = data_903 * coeffs_903;
  wire [63:0] _result_T_905 = data_904 * coeffs_904;
  wire [63:0] _result_T_906 = data_905 * coeffs_905;
  wire [63:0] _result_T_907 = data_906 * coeffs_906;
  wire [63:0] _result_T_908 = data_907 * coeffs_907;
  wire [63:0] _result_T_909 = data_908 * coeffs_908;
  wire [63:0] _result_T_910 = data_909 * coeffs_909;
  wire [63:0] _result_T_911 = data_910 * coeffs_910;
  wire [63:0] _result_T_912 = data_911 * coeffs_911;
  wire [63:0] _result_T_913 = data_912 * coeffs_912;
  wire [63:0] _result_T_914 = data_913 * coeffs_913;
  wire [63:0] _result_T_915 = data_914 * coeffs_914;
  wire [63:0] _result_T_916 = data_915 * coeffs_915;
  wire [63:0] _result_T_917 = data_916 * coeffs_916;
  wire [63:0] _result_T_918 = data_917 * coeffs_917;
  wire [63:0] _result_T_919 = data_918 * coeffs_918;
  wire [63:0] _result_T_920 = data_919 * coeffs_919;
  wire [63:0] _result_T_921 = data_920 * coeffs_920;
  wire [63:0] _result_T_922 = data_921 * coeffs_921;
  wire [63:0] _result_T_923 = data_922 * coeffs_922;
  wire [63:0] _result_T_924 = data_923 * coeffs_923;
  wire [63:0] _result_T_925 = data_924 * coeffs_924;
  wire [63:0] _result_T_926 = data_925 * coeffs_925;
  wire [63:0] _result_T_927 = data_926 * coeffs_926;
  wire [63:0] _result_T_928 = data_927 * coeffs_927;
  wire [63:0] _result_T_929 = data_928 * coeffs_928;
  wire [63:0] _result_T_930 = data_929 * coeffs_929;
  wire [63:0] _result_T_931 = data_930 * coeffs_930;
  wire [63:0] _result_T_932 = data_931 * coeffs_931;
  wire [63:0] _result_T_933 = data_932 * coeffs_932;
  wire [63:0] _result_T_934 = data_933 * coeffs_933;
  wire [63:0] _result_T_935 = data_934 * coeffs_934;
  wire [63:0] _result_T_936 = data_935 * coeffs_935;
  wire [63:0] _result_T_937 = data_936 * coeffs_936;
  wire [63:0] _result_T_938 = data_937 * coeffs_937;
  wire [63:0] _result_T_939 = data_938 * coeffs_938;
  wire [63:0] _result_T_940 = data_939 * coeffs_939;
  wire [63:0] _result_T_941 = data_940 * coeffs_940;
  wire [63:0] _result_T_942 = data_941 * coeffs_941;
  wire [63:0] _result_T_943 = data_942 * coeffs_942;
  wire [63:0] _result_T_944 = data_943 * coeffs_943;
  wire [63:0] _result_T_945 = data_944 * coeffs_944;
  wire [63:0] _result_T_946 = data_945 * coeffs_945;
  wire [63:0] _result_T_947 = data_946 * coeffs_946;
  wire [63:0] _result_T_948 = data_947 * coeffs_947;
  wire [63:0] _result_T_949 = data_948 * coeffs_948;
  wire [63:0] _result_T_950 = data_949 * coeffs_949;
  wire [63:0] _result_T_951 = data_950 * coeffs_950;
  wire [63:0] _result_T_952 = data_951 * coeffs_951;
  wire [63:0] _result_T_953 = data_952 * coeffs_952;
  wire [63:0] _result_T_954 = data_953 * coeffs_953;
  wire [63:0] _result_T_955 = data_954 * coeffs_954;
  wire [63:0] _result_T_956 = data_955 * coeffs_955;
  wire [63:0] _result_T_957 = data_956 * coeffs_956;
  wire [63:0] _result_T_958 = data_957 * coeffs_957;
  wire [63:0] _result_T_959 = data_958 * coeffs_958;
  wire [63:0] _result_T_960 = data_959 * coeffs_959;
  wire [63:0] _result_T_961 = data_960 * coeffs_960;
  wire [63:0] _result_T_962 = data_961 * coeffs_961;
  wire [63:0] _result_T_963 = data_962 * coeffs_962;
  wire [63:0] _result_T_964 = data_963 * coeffs_963;
  wire [63:0] _result_T_965 = data_964 * coeffs_964;
  wire [63:0] _result_T_966 = data_965 * coeffs_965;
  wire [63:0] _result_T_967 = data_966 * coeffs_966;
  wire [63:0] _result_T_968 = data_967 * coeffs_967;
  wire [63:0] _result_T_969 = data_968 * coeffs_968;
  wire [63:0] _result_T_970 = data_969 * coeffs_969;
  wire [63:0] _result_T_971 = data_970 * coeffs_970;
  wire [63:0] _result_T_972 = data_971 * coeffs_971;
  wire [63:0] _result_T_973 = data_972 * coeffs_972;
  wire [63:0] _result_T_974 = data_973 * coeffs_973;
  wire [63:0] _result_T_975 = data_974 * coeffs_974;
  wire [63:0] _result_T_976 = data_975 * coeffs_975;
  wire [63:0] _result_T_977 = data_976 * coeffs_976;
  wire [63:0] _result_T_978 = data_977 * coeffs_977;
  wire [63:0] _result_T_979 = data_978 * coeffs_978;
  wire [63:0] _result_T_980 = data_979 * coeffs_979;
  wire [63:0] _result_T_981 = data_980 * coeffs_980;
  wire [63:0] _result_T_982 = data_981 * coeffs_981;
  wire [63:0] _result_T_983 = data_982 * coeffs_982;
  wire [63:0] _result_T_984 = data_983 * coeffs_983;
  wire [63:0] _result_T_985 = data_984 * coeffs_984;
  wire [63:0] _result_T_986 = data_985 * coeffs_985;
  wire [63:0] _result_T_987 = data_986 * coeffs_986;
  wire [63:0] _result_T_988 = data_987 * coeffs_987;
  wire [63:0] _result_T_989 = data_988 * coeffs_988;
  wire [63:0] _result_T_990 = data_989 * coeffs_989;
  wire [63:0] _result_T_991 = data_990 * coeffs_990;
  wire [63:0] _result_T_992 = data_991 * coeffs_991;
  wire [63:0] _result_T_993 = data_992 * coeffs_992;
  wire [63:0] _result_T_994 = data_993 * coeffs_993;
  wire [63:0] _result_T_995 = data_994 * coeffs_994;
  wire [63:0] _result_T_996 = data_995 * coeffs_995;
  wire [63:0] _result_T_997 = data_996 * coeffs_996;
  wire [63:0] _result_T_998 = data_997 * coeffs_997;
  wire [63:0] _result_T_999 = data_998 * coeffs_998;
  wire [63:0] _result_T_1000 = data_999 * coeffs_999;
  wire [63:0] _result_T_1002 = _result_T_1 + _result_T_2;
  wire [63:0] _result_T_1004 = _result_T_1002 + _result_T_3;
  wire [63:0] _result_T_1006 = _result_T_1004 + _result_T_4;
  wire [63:0] _result_T_1008 = _result_T_1006 + _result_T_5;
  wire [63:0] _result_T_1010 = _result_T_1008 + _result_T_6;
  wire [63:0] _result_T_1012 = _result_T_1010 + _result_T_7;
  wire [63:0] _result_T_1014 = _result_T_1012 + _result_T_8;
  wire [63:0] _result_T_1016 = _result_T_1014 + _result_T_9;
  wire [63:0] _result_T_1018 = _result_T_1016 + _result_T_10;
  wire [63:0] _result_T_1020 = _result_T_1018 + _result_T_11;
  wire [63:0] _result_T_1022 = _result_T_1020 + _result_T_12;
  wire [63:0] _result_T_1024 = _result_T_1022 + _result_T_13;
  wire [63:0] _result_T_1026 = _result_T_1024 + _result_T_14;
  wire [63:0] _result_T_1028 = _result_T_1026 + _result_T_15;
  wire [63:0] _result_T_1030 = _result_T_1028 + _result_T_16;
  wire [63:0] _result_T_1032 = _result_T_1030 + _result_T_17;
  wire [63:0] _result_T_1034 = _result_T_1032 + _result_T_18;
  wire [63:0] _result_T_1036 = _result_T_1034 + _result_T_19;
  wire [63:0] _result_T_1038 = _result_T_1036 + _result_T_20;
  wire [63:0] _result_T_1040 = _result_T_1038 + _result_T_21;
  wire [63:0] _result_T_1042 = _result_T_1040 + _result_T_22;
  wire [63:0] _result_T_1044 = _result_T_1042 + _result_T_23;
  wire [63:0] _result_T_1046 = _result_T_1044 + _result_T_24;
  wire [63:0] _result_T_1048 = _result_T_1046 + _result_T_25;
  wire [63:0] _result_T_1050 = _result_T_1048 + _result_T_26;
  wire [63:0] _result_T_1052 = _result_T_1050 + _result_T_27;
  wire [63:0] _result_T_1054 = _result_T_1052 + _result_T_28;
  wire [63:0] _result_T_1056 = _result_T_1054 + _result_T_29;
  wire [63:0] _result_T_1058 = _result_T_1056 + _result_T_30;
  wire [63:0] _result_T_1060 = _result_T_1058 + _result_T_31;
  wire [63:0] _result_T_1062 = _result_T_1060 + _result_T_32;
  wire [63:0] _result_T_1064 = _result_T_1062 + _result_T_33;
  wire [63:0] _result_T_1066 = _result_T_1064 + _result_T_34;
  wire [63:0] _result_T_1068 = _result_T_1066 + _result_T_35;
  wire [63:0] _result_T_1070 = _result_T_1068 + _result_T_36;
  wire [63:0] _result_T_1072 = _result_T_1070 + _result_T_37;
  wire [63:0] _result_T_1074 = _result_T_1072 + _result_T_38;
  wire [63:0] _result_T_1076 = _result_T_1074 + _result_T_39;
  wire [63:0] _result_T_1078 = _result_T_1076 + _result_T_40;
  wire [63:0] _result_T_1080 = _result_T_1078 + _result_T_41;
  wire [63:0] _result_T_1082 = _result_T_1080 + _result_T_42;
  wire [63:0] _result_T_1084 = _result_T_1082 + _result_T_43;
  wire [63:0] _result_T_1086 = _result_T_1084 + _result_T_44;
  wire [63:0] _result_T_1088 = _result_T_1086 + _result_T_45;
  wire [63:0] _result_T_1090 = _result_T_1088 + _result_T_46;
  wire [63:0] _result_T_1092 = _result_T_1090 + _result_T_47;
  wire [63:0] _result_T_1094 = _result_T_1092 + _result_T_48;
  wire [63:0] _result_T_1096 = _result_T_1094 + _result_T_49;
  wire [63:0] _result_T_1098 = _result_T_1096 + _result_T_50;
  wire [63:0] _result_T_1100 = _result_T_1098 + _result_T_51;
  wire [63:0] _result_T_1102 = _result_T_1100 + _result_T_52;
  wire [63:0] _result_T_1104 = _result_T_1102 + _result_T_53;
  wire [63:0] _result_T_1106 = _result_T_1104 + _result_T_54;
  wire [63:0] _result_T_1108 = _result_T_1106 + _result_T_55;
  wire [63:0] _result_T_1110 = _result_T_1108 + _result_T_56;
  wire [63:0] _result_T_1112 = _result_T_1110 + _result_T_57;
  wire [63:0] _result_T_1114 = _result_T_1112 + _result_T_58;
  wire [63:0] _result_T_1116 = _result_T_1114 + _result_T_59;
  wire [63:0] _result_T_1118 = _result_T_1116 + _result_T_60;
  wire [63:0] _result_T_1120 = _result_T_1118 + _result_T_61;
  wire [63:0] _result_T_1122 = _result_T_1120 + _result_T_62;
  wire [63:0] _result_T_1124 = _result_T_1122 + _result_T_63;
  wire [63:0] _result_T_1126 = _result_T_1124 + _result_T_64;
  wire [63:0] _result_T_1128 = _result_T_1126 + _result_T_65;
  wire [63:0] _result_T_1130 = _result_T_1128 + _result_T_66;
  wire [63:0] _result_T_1132 = _result_T_1130 + _result_T_67;
  wire [63:0] _result_T_1134 = _result_T_1132 + _result_T_68;
  wire [63:0] _result_T_1136 = _result_T_1134 + _result_T_69;
  wire [63:0] _result_T_1138 = _result_T_1136 + _result_T_70;
  wire [63:0] _result_T_1140 = _result_T_1138 + _result_T_71;
  wire [63:0] _result_T_1142 = _result_T_1140 + _result_T_72;
  wire [63:0] _result_T_1144 = _result_T_1142 + _result_T_73;
  wire [63:0] _result_T_1146 = _result_T_1144 + _result_T_74;
  wire [63:0] _result_T_1148 = _result_T_1146 + _result_T_75;
  wire [63:0] _result_T_1150 = _result_T_1148 + _result_T_76;
  wire [63:0] _result_T_1152 = _result_T_1150 + _result_T_77;
  wire [63:0] _result_T_1154 = _result_T_1152 + _result_T_78;
  wire [63:0] _result_T_1156 = _result_T_1154 + _result_T_79;
  wire [63:0] _result_T_1158 = _result_T_1156 + _result_T_80;
  wire [63:0] _result_T_1160 = _result_T_1158 + _result_T_81;
  wire [63:0] _result_T_1162 = _result_T_1160 + _result_T_82;
  wire [63:0] _result_T_1164 = _result_T_1162 + _result_T_83;
  wire [63:0] _result_T_1166 = _result_T_1164 + _result_T_84;
  wire [63:0] _result_T_1168 = _result_T_1166 + _result_T_85;
  wire [63:0] _result_T_1170 = _result_T_1168 + _result_T_86;
  wire [63:0] _result_T_1172 = _result_T_1170 + _result_T_87;
  wire [63:0] _result_T_1174 = _result_T_1172 + _result_T_88;
  wire [63:0] _result_T_1176 = _result_T_1174 + _result_T_89;
  wire [63:0] _result_T_1178 = _result_T_1176 + _result_T_90;
  wire [63:0] _result_T_1180 = _result_T_1178 + _result_T_91;
  wire [63:0] _result_T_1182 = _result_T_1180 + _result_T_92;
  wire [63:0] _result_T_1184 = _result_T_1182 + _result_T_93;
  wire [63:0] _result_T_1186 = _result_T_1184 + _result_T_94;
  wire [63:0] _result_T_1188 = _result_T_1186 + _result_T_95;
  wire [63:0] _result_T_1190 = _result_T_1188 + _result_T_96;
  wire [63:0] _result_T_1192 = _result_T_1190 + _result_T_97;
  wire [63:0] _result_T_1194 = _result_T_1192 + _result_T_98;
  wire [63:0] _result_T_1196 = _result_T_1194 + _result_T_99;
  wire [63:0] _result_T_1198 = _result_T_1196 + _result_T_100;
  wire [63:0] _result_T_1200 = _result_T_1198 + _result_T_101;
  wire [63:0] _result_T_1202 = _result_T_1200 + _result_T_102;
  wire [63:0] _result_T_1204 = _result_T_1202 + _result_T_103;
  wire [63:0] _result_T_1206 = _result_T_1204 + _result_T_104;
  wire [63:0] _result_T_1208 = _result_T_1206 + _result_T_105;
  wire [63:0] _result_T_1210 = _result_T_1208 + _result_T_106;
  wire [63:0] _result_T_1212 = _result_T_1210 + _result_T_107;
  wire [63:0] _result_T_1214 = _result_T_1212 + _result_T_108;
  wire [63:0] _result_T_1216 = _result_T_1214 + _result_T_109;
  wire [63:0] _result_T_1218 = _result_T_1216 + _result_T_110;
  wire [63:0] _result_T_1220 = _result_T_1218 + _result_T_111;
  wire [63:0] _result_T_1222 = _result_T_1220 + _result_T_112;
  wire [63:0] _result_T_1224 = _result_T_1222 + _result_T_113;
  wire [63:0] _result_T_1226 = _result_T_1224 + _result_T_114;
  wire [63:0] _result_T_1228 = _result_T_1226 + _result_T_115;
  wire [63:0] _result_T_1230 = _result_T_1228 + _result_T_116;
  wire [63:0] _result_T_1232 = _result_T_1230 + _result_T_117;
  wire [63:0] _result_T_1234 = _result_T_1232 + _result_T_118;
  wire [63:0] _result_T_1236 = _result_T_1234 + _result_T_119;
  wire [63:0] _result_T_1238 = _result_T_1236 + _result_T_120;
  wire [63:0] _result_T_1240 = _result_T_1238 + _result_T_121;
  wire [63:0] _result_T_1242 = _result_T_1240 + _result_T_122;
  wire [63:0] _result_T_1244 = _result_T_1242 + _result_T_123;
  wire [63:0] _result_T_1246 = _result_T_1244 + _result_T_124;
  wire [63:0] _result_T_1248 = _result_T_1246 + _result_T_125;
  wire [63:0] _result_T_1250 = _result_T_1248 + _result_T_126;
  wire [63:0] _result_T_1252 = _result_T_1250 + _result_T_127;
  wire [63:0] _result_T_1254 = _result_T_1252 + _result_T_128;
  wire [63:0] _result_T_1256 = _result_T_1254 + _result_T_129;
  wire [63:0] _result_T_1258 = _result_T_1256 + _result_T_130;
  wire [63:0] _result_T_1260 = _result_T_1258 + _result_T_131;
  wire [63:0] _result_T_1262 = _result_T_1260 + _result_T_132;
  wire [63:0] _result_T_1264 = _result_T_1262 + _result_T_133;
  wire [63:0] _result_T_1266 = _result_T_1264 + _result_T_134;
  wire [63:0] _result_T_1268 = _result_T_1266 + _result_T_135;
  wire [63:0] _result_T_1270 = _result_T_1268 + _result_T_136;
  wire [63:0] _result_T_1272 = _result_T_1270 + _result_T_137;
  wire [63:0] _result_T_1274 = _result_T_1272 + _result_T_138;
  wire [63:0] _result_T_1276 = _result_T_1274 + _result_T_139;
  wire [63:0] _result_T_1278 = _result_T_1276 + _result_T_140;
  wire [63:0] _result_T_1280 = _result_T_1278 + _result_T_141;
  wire [63:0] _result_T_1282 = _result_T_1280 + _result_T_142;
  wire [63:0] _result_T_1284 = _result_T_1282 + _result_T_143;
  wire [63:0] _result_T_1286 = _result_T_1284 + _result_T_144;
  wire [63:0] _result_T_1288 = _result_T_1286 + _result_T_145;
  wire [63:0] _result_T_1290 = _result_T_1288 + _result_T_146;
  wire [63:0] _result_T_1292 = _result_T_1290 + _result_T_147;
  wire [63:0] _result_T_1294 = _result_T_1292 + _result_T_148;
  wire [63:0] _result_T_1296 = _result_T_1294 + _result_T_149;
  wire [63:0] _result_T_1298 = _result_T_1296 + _result_T_150;
  wire [63:0] _result_T_1300 = _result_T_1298 + _result_T_151;
  wire [63:0] _result_T_1302 = _result_T_1300 + _result_T_152;
  wire [63:0] _result_T_1304 = _result_T_1302 + _result_T_153;
  wire [63:0] _result_T_1306 = _result_T_1304 + _result_T_154;
  wire [63:0] _result_T_1308 = _result_T_1306 + _result_T_155;
  wire [63:0] _result_T_1310 = _result_T_1308 + _result_T_156;
  wire [63:0] _result_T_1312 = _result_T_1310 + _result_T_157;
  wire [63:0] _result_T_1314 = _result_T_1312 + _result_T_158;
  wire [63:0] _result_T_1316 = _result_T_1314 + _result_T_159;
  wire [63:0] _result_T_1318 = _result_T_1316 + _result_T_160;
  wire [63:0] _result_T_1320 = _result_T_1318 + _result_T_161;
  wire [63:0] _result_T_1322 = _result_T_1320 + _result_T_162;
  wire [63:0] _result_T_1324 = _result_T_1322 + _result_T_163;
  wire [63:0] _result_T_1326 = _result_T_1324 + _result_T_164;
  wire [63:0] _result_T_1328 = _result_T_1326 + _result_T_165;
  wire [63:0] _result_T_1330 = _result_T_1328 + _result_T_166;
  wire [63:0] _result_T_1332 = _result_T_1330 + _result_T_167;
  wire [63:0] _result_T_1334 = _result_T_1332 + _result_T_168;
  wire [63:0] _result_T_1336 = _result_T_1334 + _result_T_169;
  wire [63:0] _result_T_1338 = _result_T_1336 + _result_T_170;
  wire [63:0] _result_T_1340 = _result_T_1338 + _result_T_171;
  wire [63:0] _result_T_1342 = _result_T_1340 + _result_T_172;
  wire [63:0] _result_T_1344 = _result_T_1342 + _result_T_173;
  wire [63:0] _result_T_1346 = _result_T_1344 + _result_T_174;
  wire [63:0] _result_T_1348 = _result_T_1346 + _result_T_175;
  wire [63:0] _result_T_1350 = _result_T_1348 + _result_T_176;
  wire [63:0] _result_T_1352 = _result_T_1350 + _result_T_177;
  wire [63:0] _result_T_1354 = _result_T_1352 + _result_T_178;
  wire [63:0] _result_T_1356 = _result_T_1354 + _result_T_179;
  wire [63:0] _result_T_1358 = _result_T_1356 + _result_T_180;
  wire [63:0] _result_T_1360 = _result_T_1358 + _result_T_181;
  wire [63:0] _result_T_1362 = _result_T_1360 + _result_T_182;
  wire [63:0] _result_T_1364 = _result_T_1362 + _result_T_183;
  wire [63:0] _result_T_1366 = _result_T_1364 + _result_T_184;
  wire [63:0] _result_T_1368 = _result_T_1366 + _result_T_185;
  wire [63:0] _result_T_1370 = _result_T_1368 + _result_T_186;
  wire [63:0] _result_T_1372 = _result_T_1370 + _result_T_187;
  wire [63:0] _result_T_1374 = _result_T_1372 + _result_T_188;
  wire [63:0] _result_T_1376 = _result_T_1374 + _result_T_189;
  wire [63:0] _result_T_1378 = _result_T_1376 + _result_T_190;
  wire [63:0] _result_T_1380 = _result_T_1378 + _result_T_191;
  wire [63:0] _result_T_1382 = _result_T_1380 + _result_T_192;
  wire [63:0] _result_T_1384 = _result_T_1382 + _result_T_193;
  wire [63:0] _result_T_1386 = _result_T_1384 + _result_T_194;
  wire [63:0] _result_T_1388 = _result_T_1386 + _result_T_195;
  wire [63:0] _result_T_1390 = _result_T_1388 + _result_T_196;
  wire [63:0] _result_T_1392 = _result_T_1390 + _result_T_197;
  wire [63:0] _result_T_1394 = _result_T_1392 + _result_T_198;
  wire [63:0] _result_T_1396 = _result_T_1394 + _result_T_199;
  wire [63:0] _result_T_1398 = _result_T_1396 + _result_T_200;
  wire [63:0] _result_T_1400 = _result_T_1398 + _result_T_201;
  wire [63:0] _result_T_1402 = _result_T_1400 + _result_T_202;
  wire [63:0] _result_T_1404 = _result_T_1402 + _result_T_203;
  wire [63:0] _result_T_1406 = _result_T_1404 + _result_T_204;
  wire [63:0] _result_T_1408 = _result_T_1406 + _result_T_205;
  wire [63:0] _result_T_1410 = _result_T_1408 + _result_T_206;
  wire [63:0] _result_T_1412 = _result_T_1410 + _result_T_207;
  wire [63:0] _result_T_1414 = _result_T_1412 + _result_T_208;
  wire [63:0] _result_T_1416 = _result_T_1414 + _result_T_209;
  wire [63:0] _result_T_1418 = _result_T_1416 + _result_T_210;
  wire [63:0] _result_T_1420 = _result_T_1418 + _result_T_211;
  wire [63:0] _result_T_1422 = _result_T_1420 + _result_T_212;
  wire [63:0] _result_T_1424 = _result_T_1422 + _result_T_213;
  wire [63:0] _result_T_1426 = _result_T_1424 + _result_T_214;
  wire [63:0] _result_T_1428 = _result_T_1426 + _result_T_215;
  wire [63:0] _result_T_1430 = _result_T_1428 + _result_T_216;
  wire [63:0] _result_T_1432 = _result_T_1430 + _result_T_217;
  wire [63:0] _result_T_1434 = _result_T_1432 + _result_T_218;
  wire [63:0] _result_T_1436 = _result_T_1434 + _result_T_219;
  wire [63:0] _result_T_1438 = _result_T_1436 + _result_T_220;
  wire [63:0] _result_T_1440 = _result_T_1438 + _result_T_221;
  wire [63:0] _result_T_1442 = _result_T_1440 + _result_T_222;
  wire [63:0] _result_T_1444 = _result_T_1442 + _result_T_223;
  wire [63:0] _result_T_1446 = _result_T_1444 + _result_T_224;
  wire [63:0] _result_T_1448 = _result_T_1446 + _result_T_225;
  wire [63:0] _result_T_1450 = _result_T_1448 + _result_T_226;
  wire [63:0] _result_T_1452 = _result_T_1450 + _result_T_227;
  wire [63:0] _result_T_1454 = _result_T_1452 + _result_T_228;
  wire [63:0] _result_T_1456 = _result_T_1454 + _result_T_229;
  wire [63:0] _result_T_1458 = _result_T_1456 + _result_T_230;
  wire [63:0] _result_T_1460 = _result_T_1458 + _result_T_231;
  wire [63:0] _result_T_1462 = _result_T_1460 + _result_T_232;
  wire [63:0] _result_T_1464 = _result_T_1462 + _result_T_233;
  wire [63:0] _result_T_1466 = _result_T_1464 + _result_T_234;
  wire [63:0] _result_T_1468 = _result_T_1466 + _result_T_235;
  wire [63:0] _result_T_1470 = _result_T_1468 + _result_T_236;
  wire [63:0] _result_T_1472 = _result_T_1470 + _result_T_237;
  wire [63:0] _result_T_1474 = _result_T_1472 + _result_T_238;
  wire [63:0] _result_T_1476 = _result_T_1474 + _result_T_239;
  wire [63:0] _result_T_1478 = _result_T_1476 + _result_T_240;
  wire [63:0] _result_T_1480 = _result_T_1478 + _result_T_241;
  wire [63:0] _result_T_1482 = _result_T_1480 + _result_T_242;
  wire [63:0] _result_T_1484 = _result_T_1482 + _result_T_243;
  wire [63:0] _result_T_1486 = _result_T_1484 + _result_T_244;
  wire [63:0] _result_T_1488 = _result_T_1486 + _result_T_245;
  wire [63:0] _result_T_1490 = _result_T_1488 + _result_T_246;
  wire [63:0] _result_T_1492 = _result_T_1490 + _result_T_247;
  wire [63:0] _result_T_1494 = _result_T_1492 + _result_T_248;
  wire [63:0] _result_T_1496 = _result_T_1494 + _result_T_249;
  wire [63:0] _result_T_1498 = _result_T_1496 + _result_T_250;
  wire [63:0] _result_T_1500 = _result_T_1498 + _result_T_251;
  wire [63:0] _result_T_1502 = _result_T_1500 + _result_T_252;
  wire [63:0] _result_T_1504 = _result_T_1502 + _result_T_253;
  wire [63:0] _result_T_1506 = _result_T_1504 + _result_T_254;
  wire [63:0] _result_T_1508 = _result_T_1506 + _result_T_255;
  wire [63:0] _result_T_1510 = _result_T_1508 + _result_T_256;
  wire [63:0] _result_T_1512 = _result_T_1510 + _result_T_257;
  wire [63:0] _result_T_1514 = _result_T_1512 + _result_T_258;
  wire [63:0] _result_T_1516 = _result_T_1514 + _result_T_259;
  wire [63:0] _result_T_1518 = _result_T_1516 + _result_T_260;
  wire [63:0] _result_T_1520 = _result_T_1518 + _result_T_261;
  wire [63:0] _result_T_1522 = _result_T_1520 + _result_T_262;
  wire [63:0] _result_T_1524 = _result_T_1522 + _result_T_263;
  wire [63:0] _result_T_1526 = _result_T_1524 + _result_T_264;
  wire [63:0] _result_T_1528 = _result_T_1526 + _result_T_265;
  wire [63:0] _result_T_1530 = _result_T_1528 + _result_T_266;
  wire [63:0] _result_T_1532 = _result_T_1530 + _result_T_267;
  wire [63:0] _result_T_1534 = _result_T_1532 + _result_T_268;
  wire [63:0] _result_T_1536 = _result_T_1534 + _result_T_269;
  wire [63:0] _result_T_1538 = _result_T_1536 + _result_T_270;
  wire [63:0] _result_T_1540 = _result_T_1538 + _result_T_271;
  wire [63:0] _result_T_1542 = _result_T_1540 + _result_T_272;
  wire [63:0] _result_T_1544 = _result_T_1542 + _result_T_273;
  wire [63:0] _result_T_1546 = _result_T_1544 + _result_T_274;
  wire [63:0] _result_T_1548 = _result_T_1546 + _result_T_275;
  wire [63:0] _result_T_1550 = _result_T_1548 + _result_T_276;
  wire [63:0] _result_T_1552 = _result_T_1550 + _result_T_277;
  wire [63:0] _result_T_1554 = _result_T_1552 + _result_T_278;
  wire [63:0] _result_T_1556 = _result_T_1554 + _result_T_279;
  wire [63:0] _result_T_1558 = _result_T_1556 + _result_T_280;
  wire [63:0] _result_T_1560 = _result_T_1558 + _result_T_281;
  wire [63:0] _result_T_1562 = _result_T_1560 + _result_T_282;
  wire [63:0] _result_T_1564 = _result_T_1562 + _result_T_283;
  wire [63:0] _result_T_1566 = _result_T_1564 + _result_T_284;
  wire [63:0] _result_T_1568 = _result_T_1566 + _result_T_285;
  wire [63:0] _result_T_1570 = _result_T_1568 + _result_T_286;
  wire [63:0] _result_T_1572 = _result_T_1570 + _result_T_287;
  wire [63:0] _result_T_1574 = _result_T_1572 + _result_T_288;
  wire [63:0] _result_T_1576 = _result_T_1574 + _result_T_289;
  wire [63:0] _result_T_1578 = _result_T_1576 + _result_T_290;
  wire [63:0] _result_T_1580 = _result_T_1578 + _result_T_291;
  wire [63:0] _result_T_1582 = _result_T_1580 + _result_T_292;
  wire [63:0] _result_T_1584 = _result_T_1582 + _result_T_293;
  wire [63:0] _result_T_1586 = _result_T_1584 + _result_T_294;
  wire [63:0] _result_T_1588 = _result_T_1586 + _result_T_295;
  wire [63:0] _result_T_1590 = _result_T_1588 + _result_T_296;
  wire [63:0] _result_T_1592 = _result_T_1590 + _result_T_297;
  wire [63:0] _result_T_1594 = _result_T_1592 + _result_T_298;
  wire [63:0] _result_T_1596 = _result_T_1594 + _result_T_299;
  wire [63:0] _result_T_1598 = _result_T_1596 + _result_T_300;
  wire [63:0] _result_T_1600 = _result_T_1598 + _result_T_301;
  wire [63:0] _result_T_1602 = _result_T_1600 + _result_T_302;
  wire [63:0] _result_T_1604 = _result_T_1602 + _result_T_303;
  wire [63:0] _result_T_1606 = _result_T_1604 + _result_T_304;
  wire [63:0] _result_T_1608 = _result_T_1606 + _result_T_305;
  wire [63:0] _result_T_1610 = _result_T_1608 + _result_T_306;
  wire [63:0] _result_T_1612 = _result_T_1610 + _result_T_307;
  wire [63:0] _result_T_1614 = _result_T_1612 + _result_T_308;
  wire [63:0] _result_T_1616 = _result_T_1614 + _result_T_309;
  wire [63:0] _result_T_1618 = _result_T_1616 + _result_T_310;
  wire [63:0] _result_T_1620 = _result_T_1618 + _result_T_311;
  wire [63:0] _result_T_1622 = _result_T_1620 + _result_T_312;
  wire [63:0] _result_T_1624 = _result_T_1622 + _result_T_313;
  wire [63:0] _result_T_1626 = _result_T_1624 + _result_T_314;
  wire [63:0] _result_T_1628 = _result_T_1626 + _result_T_315;
  wire [63:0] _result_T_1630 = _result_T_1628 + _result_T_316;
  wire [63:0] _result_T_1632 = _result_T_1630 + _result_T_317;
  wire [63:0] _result_T_1634 = _result_T_1632 + _result_T_318;
  wire [63:0] _result_T_1636 = _result_T_1634 + _result_T_319;
  wire [63:0] _result_T_1638 = _result_T_1636 + _result_T_320;
  wire [63:0] _result_T_1640 = _result_T_1638 + _result_T_321;
  wire [63:0] _result_T_1642 = _result_T_1640 + _result_T_322;
  wire [63:0] _result_T_1644 = _result_T_1642 + _result_T_323;
  wire [63:0] _result_T_1646 = _result_T_1644 + _result_T_324;
  wire [63:0] _result_T_1648 = _result_T_1646 + _result_T_325;
  wire [63:0] _result_T_1650 = _result_T_1648 + _result_T_326;
  wire [63:0] _result_T_1652 = _result_T_1650 + _result_T_327;
  wire [63:0] _result_T_1654 = _result_T_1652 + _result_T_328;
  wire [63:0] _result_T_1656 = _result_T_1654 + _result_T_329;
  wire [63:0] _result_T_1658 = _result_T_1656 + _result_T_330;
  wire [63:0] _result_T_1660 = _result_T_1658 + _result_T_331;
  wire [63:0] _result_T_1662 = _result_T_1660 + _result_T_332;
  wire [63:0] _result_T_1664 = _result_T_1662 + _result_T_333;
  wire [63:0] _result_T_1666 = _result_T_1664 + _result_T_334;
  wire [63:0] _result_T_1668 = _result_T_1666 + _result_T_335;
  wire [63:0] _result_T_1670 = _result_T_1668 + _result_T_336;
  wire [63:0] _result_T_1672 = _result_T_1670 + _result_T_337;
  wire [63:0] _result_T_1674 = _result_T_1672 + _result_T_338;
  wire [63:0] _result_T_1676 = _result_T_1674 + _result_T_339;
  wire [63:0] _result_T_1678 = _result_T_1676 + _result_T_340;
  wire [63:0] _result_T_1680 = _result_T_1678 + _result_T_341;
  wire [63:0] _result_T_1682 = _result_T_1680 + _result_T_342;
  wire [63:0] _result_T_1684 = _result_T_1682 + _result_T_343;
  wire [63:0] _result_T_1686 = _result_T_1684 + _result_T_344;
  wire [63:0] _result_T_1688 = _result_T_1686 + _result_T_345;
  wire [63:0] _result_T_1690 = _result_T_1688 + _result_T_346;
  wire [63:0] _result_T_1692 = _result_T_1690 + _result_T_347;
  wire [63:0] _result_T_1694 = _result_T_1692 + _result_T_348;
  wire [63:0] _result_T_1696 = _result_T_1694 + _result_T_349;
  wire [63:0] _result_T_1698 = _result_T_1696 + _result_T_350;
  wire [63:0] _result_T_1700 = _result_T_1698 + _result_T_351;
  wire [63:0] _result_T_1702 = _result_T_1700 + _result_T_352;
  wire [63:0] _result_T_1704 = _result_T_1702 + _result_T_353;
  wire [63:0] _result_T_1706 = _result_T_1704 + _result_T_354;
  wire [63:0] _result_T_1708 = _result_T_1706 + _result_T_355;
  wire [63:0] _result_T_1710 = _result_T_1708 + _result_T_356;
  wire [63:0] _result_T_1712 = _result_T_1710 + _result_T_357;
  wire [63:0] _result_T_1714 = _result_T_1712 + _result_T_358;
  wire [63:0] _result_T_1716 = _result_T_1714 + _result_T_359;
  wire [63:0] _result_T_1718 = _result_T_1716 + _result_T_360;
  wire [63:0] _result_T_1720 = _result_T_1718 + _result_T_361;
  wire [63:0] _result_T_1722 = _result_T_1720 + _result_T_362;
  wire [63:0] _result_T_1724 = _result_T_1722 + _result_T_363;
  wire [63:0] _result_T_1726 = _result_T_1724 + _result_T_364;
  wire [63:0] _result_T_1728 = _result_T_1726 + _result_T_365;
  wire [63:0] _result_T_1730 = _result_T_1728 + _result_T_366;
  wire [63:0] _result_T_1732 = _result_T_1730 + _result_T_367;
  wire [63:0] _result_T_1734 = _result_T_1732 + _result_T_368;
  wire [63:0] _result_T_1736 = _result_T_1734 + _result_T_369;
  wire [63:0] _result_T_1738 = _result_T_1736 + _result_T_370;
  wire [63:0] _result_T_1740 = _result_T_1738 + _result_T_371;
  wire [63:0] _result_T_1742 = _result_T_1740 + _result_T_372;
  wire [63:0] _result_T_1744 = _result_T_1742 + _result_T_373;
  wire [63:0] _result_T_1746 = _result_T_1744 + _result_T_374;
  wire [63:0] _result_T_1748 = _result_T_1746 + _result_T_375;
  wire [63:0] _result_T_1750 = _result_T_1748 + _result_T_376;
  wire [63:0] _result_T_1752 = _result_T_1750 + _result_T_377;
  wire [63:0] _result_T_1754 = _result_T_1752 + _result_T_378;
  wire [63:0] _result_T_1756 = _result_T_1754 + _result_T_379;
  wire [63:0] _result_T_1758 = _result_T_1756 + _result_T_380;
  wire [63:0] _result_T_1760 = _result_T_1758 + _result_T_381;
  wire [63:0] _result_T_1762 = _result_T_1760 + _result_T_382;
  wire [63:0] _result_T_1764 = _result_T_1762 + _result_T_383;
  wire [63:0] _result_T_1766 = _result_T_1764 + _result_T_384;
  wire [63:0] _result_T_1768 = _result_T_1766 + _result_T_385;
  wire [63:0] _result_T_1770 = _result_T_1768 + _result_T_386;
  wire [63:0] _result_T_1772 = _result_T_1770 + _result_T_387;
  wire [63:0] _result_T_1774 = _result_T_1772 + _result_T_388;
  wire [63:0] _result_T_1776 = _result_T_1774 + _result_T_389;
  wire [63:0] _result_T_1778 = _result_T_1776 + _result_T_390;
  wire [63:0] _result_T_1780 = _result_T_1778 + _result_T_391;
  wire [63:0] _result_T_1782 = _result_T_1780 + _result_T_392;
  wire [63:0] _result_T_1784 = _result_T_1782 + _result_T_393;
  wire [63:0] _result_T_1786 = _result_T_1784 + _result_T_394;
  wire [63:0] _result_T_1788 = _result_T_1786 + _result_T_395;
  wire [63:0] _result_T_1790 = _result_T_1788 + _result_T_396;
  wire [63:0] _result_T_1792 = _result_T_1790 + _result_T_397;
  wire [63:0] _result_T_1794 = _result_T_1792 + _result_T_398;
  wire [63:0] _result_T_1796 = _result_T_1794 + _result_T_399;
  wire [63:0] _result_T_1798 = _result_T_1796 + _result_T_400;
  wire [63:0] _result_T_1800 = _result_T_1798 + _result_T_401;
  wire [63:0] _result_T_1802 = _result_T_1800 + _result_T_402;
  wire [63:0] _result_T_1804 = _result_T_1802 + _result_T_403;
  wire [63:0] _result_T_1806 = _result_T_1804 + _result_T_404;
  wire [63:0] _result_T_1808 = _result_T_1806 + _result_T_405;
  wire [63:0] _result_T_1810 = _result_T_1808 + _result_T_406;
  wire [63:0] _result_T_1812 = _result_T_1810 + _result_T_407;
  wire [63:0] _result_T_1814 = _result_T_1812 + _result_T_408;
  wire [63:0] _result_T_1816 = _result_T_1814 + _result_T_409;
  wire [63:0] _result_T_1818 = _result_T_1816 + _result_T_410;
  wire [63:0] _result_T_1820 = _result_T_1818 + _result_T_411;
  wire [63:0] _result_T_1822 = _result_T_1820 + _result_T_412;
  wire [63:0] _result_T_1824 = _result_T_1822 + _result_T_413;
  wire [63:0] _result_T_1826 = _result_T_1824 + _result_T_414;
  wire [63:0] _result_T_1828 = _result_T_1826 + _result_T_415;
  wire [63:0] _result_T_1830 = _result_T_1828 + _result_T_416;
  wire [63:0] _result_T_1832 = _result_T_1830 + _result_T_417;
  wire [63:0] _result_T_1834 = _result_T_1832 + _result_T_418;
  wire [63:0] _result_T_1836 = _result_T_1834 + _result_T_419;
  wire [63:0] _result_T_1838 = _result_T_1836 + _result_T_420;
  wire [63:0] _result_T_1840 = _result_T_1838 + _result_T_421;
  wire [63:0] _result_T_1842 = _result_T_1840 + _result_T_422;
  wire [63:0] _result_T_1844 = _result_T_1842 + _result_T_423;
  wire [63:0] _result_T_1846 = _result_T_1844 + _result_T_424;
  wire [63:0] _result_T_1848 = _result_T_1846 + _result_T_425;
  wire [63:0] _result_T_1850 = _result_T_1848 + _result_T_426;
  wire [63:0] _result_T_1852 = _result_T_1850 + _result_T_427;
  wire [63:0] _result_T_1854 = _result_T_1852 + _result_T_428;
  wire [63:0] _result_T_1856 = _result_T_1854 + _result_T_429;
  wire [63:0] _result_T_1858 = _result_T_1856 + _result_T_430;
  wire [63:0] _result_T_1860 = _result_T_1858 + _result_T_431;
  wire [63:0] _result_T_1862 = _result_T_1860 + _result_T_432;
  wire [63:0] _result_T_1864 = _result_T_1862 + _result_T_433;
  wire [63:0] _result_T_1866 = _result_T_1864 + _result_T_434;
  wire [63:0] _result_T_1868 = _result_T_1866 + _result_T_435;
  wire [63:0] _result_T_1870 = _result_T_1868 + _result_T_436;
  wire [63:0] _result_T_1872 = _result_T_1870 + _result_T_437;
  wire [63:0] _result_T_1874 = _result_T_1872 + _result_T_438;
  wire [63:0] _result_T_1876 = _result_T_1874 + _result_T_439;
  wire [63:0] _result_T_1878 = _result_T_1876 + _result_T_440;
  wire [63:0] _result_T_1880 = _result_T_1878 + _result_T_441;
  wire [63:0] _result_T_1882 = _result_T_1880 + _result_T_442;
  wire [63:0] _result_T_1884 = _result_T_1882 + _result_T_443;
  wire [63:0] _result_T_1886 = _result_T_1884 + _result_T_444;
  wire [63:0] _result_T_1888 = _result_T_1886 + _result_T_445;
  wire [63:0] _result_T_1890 = _result_T_1888 + _result_T_446;
  wire [63:0] _result_T_1892 = _result_T_1890 + _result_T_447;
  wire [63:0] _result_T_1894 = _result_T_1892 + _result_T_448;
  wire [63:0] _result_T_1896 = _result_T_1894 + _result_T_449;
  wire [63:0] _result_T_1898 = _result_T_1896 + _result_T_450;
  wire [63:0] _result_T_1900 = _result_T_1898 + _result_T_451;
  wire [63:0] _result_T_1902 = _result_T_1900 + _result_T_452;
  wire [63:0] _result_T_1904 = _result_T_1902 + _result_T_453;
  wire [63:0] _result_T_1906 = _result_T_1904 + _result_T_454;
  wire [63:0] _result_T_1908 = _result_T_1906 + _result_T_455;
  wire [63:0] _result_T_1910 = _result_T_1908 + _result_T_456;
  wire [63:0] _result_T_1912 = _result_T_1910 + _result_T_457;
  wire [63:0] _result_T_1914 = _result_T_1912 + _result_T_458;
  wire [63:0] _result_T_1916 = _result_T_1914 + _result_T_459;
  wire [63:0] _result_T_1918 = _result_T_1916 + _result_T_460;
  wire [63:0] _result_T_1920 = _result_T_1918 + _result_T_461;
  wire [63:0] _result_T_1922 = _result_T_1920 + _result_T_462;
  wire [63:0] _result_T_1924 = _result_T_1922 + _result_T_463;
  wire [63:0] _result_T_1926 = _result_T_1924 + _result_T_464;
  wire [63:0] _result_T_1928 = _result_T_1926 + _result_T_465;
  wire [63:0] _result_T_1930 = _result_T_1928 + _result_T_466;
  wire [63:0] _result_T_1932 = _result_T_1930 + _result_T_467;
  wire [63:0] _result_T_1934 = _result_T_1932 + _result_T_468;
  wire [63:0] _result_T_1936 = _result_T_1934 + _result_T_469;
  wire [63:0] _result_T_1938 = _result_T_1936 + _result_T_470;
  wire [63:0] _result_T_1940 = _result_T_1938 + _result_T_471;
  wire [63:0] _result_T_1942 = _result_T_1940 + _result_T_472;
  wire [63:0] _result_T_1944 = _result_T_1942 + _result_T_473;
  wire [63:0] _result_T_1946 = _result_T_1944 + _result_T_474;
  wire [63:0] _result_T_1948 = _result_T_1946 + _result_T_475;
  wire [63:0] _result_T_1950 = _result_T_1948 + _result_T_476;
  wire [63:0] _result_T_1952 = _result_T_1950 + _result_T_477;
  wire [63:0] _result_T_1954 = _result_T_1952 + _result_T_478;
  wire [63:0] _result_T_1956 = _result_T_1954 + _result_T_479;
  wire [63:0] _result_T_1958 = _result_T_1956 + _result_T_480;
  wire [63:0] _result_T_1960 = _result_T_1958 + _result_T_481;
  wire [63:0] _result_T_1962 = _result_T_1960 + _result_T_482;
  wire [63:0] _result_T_1964 = _result_T_1962 + _result_T_483;
  wire [63:0] _result_T_1966 = _result_T_1964 + _result_T_484;
  wire [63:0] _result_T_1968 = _result_T_1966 + _result_T_485;
  wire [63:0] _result_T_1970 = _result_T_1968 + _result_T_486;
  wire [63:0] _result_T_1972 = _result_T_1970 + _result_T_487;
  wire [63:0] _result_T_1974 = _result_T_1972 + _result_T_488;
  wire [63:0] _result_T_1976 = _result_T_1974 + _result_T_489;
  wire [63:0] _result_T_1978 = _result_T_1976 + _result_T_490;
  wire [63:0] _result_T_1980 = _result_T_1978 + _result_T_491;
  wire [63:0] _result_T_1982 = _result_T_1980 + _result_T_492;
  wire [63:0] _result_T_1984 = _result_T_1982 + _result_T_493;
  wire [63:0] _result_T_1986 = _result_T_1984 + _result_T_494;
  wire [63:0] _result_T_1988 = _result_T_1986 + _result_T_495;
  wire [63:0] _result_T_1990 = _result_T_1988 + _result_T_496;
  wire [63:0] _result_T_1992 = _result_T_1990 + _result_T_497;
  wire [63:0] _result_T_1994 = _result_T_1992 + _result_T_498;
  wire [63:0] _result_T_1996 = _result_T_1994 + _result_T_499;
  wire [63:0] _result_T_1998 = _result_T_1996 + _result_T_500;
  wire [63:0] _result_T_2000 = _result_T_1998 + _result_T_501;
  wire [63:0] _result_T_2002 = _result_T_2000 + _result_T_502;
  wire [63:0] _result_T_2004 = _result_T_2002 + _result_T_503;
  wire [63:0] _result_T_2006 = _result_T_2004 + _result_T_504;
  wire [63:0] _result_T_2008 = _result_T_2006 + _result_T_505;
  wire [63:0] _result_T_2010 = _result_T_2008 + _result_T_506;
  wire [63:0] _result_T_2012 = _result_T_2010 + _result_T_507;
  wire [63:0] _result_T_2014 = _result_T_2012 + _result_T_508;
  wire [63:0] _result_T_2016 = _result_T_2014 + _result_T_509;
  wire [63:0] _result_T_2018 = _result_T_2016 + _result_T_510;
  wire [63:0] _result_T_2020 = _result_T_2018 + _result_T_511;
  wire [63:0] _result_T_2022 = _result_T_2020 + _result_T_512;
  wire [63:0] _result_T_2024 = _result_T_2022 + _result_T_513;
  wire [63:0] _result_T_2026 = _result_T_2024 + _result_T_514;
  wire [63:0] _result_T_2028 = _result_T_2026 + _result_T_515;
  wire [63:0] _result_T_2030 = _result_T_2028 + _result_T_516;
  wire [63:0] _result_T_2032 = _result_T_2030 + _result_T_517;
  wire [63:0] _result_T_2034 = _result_T_2032 + _result_T_518;
  wire [63:0] _result_T_2036 = _result_T_2034 + _result_T_519;
  wire [63:0] _result_T_2038 = _result_T_2036 + _result_T_520;
  wire [63:0] _result_T_2040 = _result_T_2038 + _result_T_521;
  wire [63:0] _result_T_2042 = _result_T_2040 + _result_T_522;
  wire [63:0] _result_T_2044 = _result_T_2042 + _result_T_523;
  wire [63:0] _result_T_2046 = _result_T_2044 + _result_T_524;
  wire [63:0] _result_T_2048 = _result_T_2046 + _result_T_525;
  wire [63:0] _result_T_2050 = _result_T_2048 + _result_T_526;
  wire [63:0] _result_T_2052 = _result_T_2050 + _result_T_527;
  wire [63:0] _result_T_2054 = _result_T_2052 + _result_T_528;
  wire [63:0] _result_T_2056 = _result_T_2054 + _result_T_529;
  wire [63:0] _result_T_2058 = _result_T_2056 + _result_T_530;
  wire [63:0] _result_T_2060 = _result_T_2058 + _result_T_531;
  wire [63:0] _result_T_2062 = _result_T_2060 + _result_T_532;
  wire [63:0] _result_T_2064 = _result_T_2062 + _result_T_533;
  wire [63:0] _result_T_2066 = _result_T_2064 + _result_T_534;
  wire [63:0] _result_T_2068 = _result_T_2066 + _result_T_535;
  wire [63:0] _result_T_2070 = _result_T_2068 + _result_T_536;
  wire [63:0] _result_T_2072 = _result_T_2070 + _result_T_537;
  wire [63:0] _result_T_2074 = _result_T_2072 + _result_T_538;
  wire [63:0] _result_T_2076 = _result_T_2074 + _result_T_539;
  wire [63:0] _result_T_2078 = _result_T_2076 + _result_T_540;
  wire [63:0] _result_T_2080 = _result_T_2078 + _result_T_541;
  wire [63:0] _result_T_2082 = _result_T_2080 + _result_T_542;
  wire [63:0] _result_T_2084 = _result_T_2082 + _result_T_543;
  wire [63:0] _result_T_2086 = _result_T_2084 + _result_T_544;
  wire [63:0] _result_T_2088 = _result_T_2086 + _result_T_545;
  wire [63:0] _result_T_2090 = _result_T_2088 + _result_T_546;
  wire [63:0] _result_T_2092 = _result_T_2090 + _result_T_547;
  wire [63:0] _result_T_2094 = _result_T_2092 + _result_T_548;
  wire [63:0] _result_T_2096 = _result_T_2094 + _result_T_549;
  wire [63:0] _result_T_2098 = _result_T_2096 + _result_T_550;
  wire [63:0] _result_T_2100 = _result_T_2098 + _result_T_551;
  wire [63:0] _result_T_2102 = _result_T_2100 + _result_T_552;
  wire [63:0] _result_T_2104 = _result_T_2102 + _result_T_553;
  wire [63:0] _result_T_2106 = _result_T_2104 + _result_T_554;
  wire [63:0] _result_T_2108 = _result_T_2106 + _result_T_555;
  wire [63:0] _result_T_2110 = _result_T_2108 + _result_T_556;
  wire [63:0] _result_T_2112 = _result_T_2110 + _result_T_557;
  wire [63:0] _result_T_2114 = _result_T_2112 + _result_T_558;
  wire [63:0] _result_T_2116 = _result_T_2114 + _result_T_559;
  wire [63:0] _result_T_2118 = _result_T_2116 + _result_T_560;
  wire [63:0] _result_T_2120 = _result_T_2118 + _result_T_561;
  wire [63:0] _result_T_2122 = _result_T_2120 + _result_T_562;
  wire [63:0] _result_T_2124 = _result_T_2122 + _result_T_563;
  wire [63:0] _result_T_2126 = _result_T_2124 + _result_T_564;
  wire [63:0] _result_T_2128 = _result_T_2126 + _result_T_565;
  wire [63:0] _result_T_2130 = _result_T_2128 + _result_T_566;
  wire [63:0] _result_T_2132 = _result_T_2130 + _result_T_567;
  wire [63:0] _result_T_2134 = _result_T_2132 + _result_T_568;
  wire [63:0] _result_T_2136 = _result_T_2134 + _result_T_569;
  wire [63:0] _result_T_2138 = _result_T_2136 + _result_T_570;
  wire [63:0] _result_T_2140 = _result_T_2138 + _result_T_571;
  wire [63:0] _result_T_2142 = _result_T_2140 + _result_T_572;
  wire [63:0] _result_T_2144 = _result_T_2142 + _result_T_573;
  wire [63:0] _result_T_2146 = _result_T_2144 + _result_T_574;
  wire [63:0] _result_T_2148 = _result_T_2146 + _result_T_575;
  wire [63:0] _result_T_2150 = _result_T_2148 + _result_T_576;
  wire [63:0] _result_T_2152 = _result_T_2150 + _result_T_577;
  wire [63:0] _result_T_2154 = _result_T_2152 + _result_T_578;
  wire [63:0] _result_T_2156 = _result_T_2154 + _result_T_579;
  wire [63:0] _result_T_2158 = _result_T_2156 + _result_T_580;
  wire [63:0] _result_T_2160 = _result_T_2158 + _result_T_581;
  wire [63:0] _result_T_2162 = _result_T_2160 + _result_T_582;
  wire [63:0] _result_T_2164 = _result_T_2162 + _result_T_583;
  wire [63:0] _result_T_2166 = _result_T_2164 + _result_T_584;
  wire [63:0] _result_T_2168 = _result_T_2166 + _result_T_585;
  wire [63:0] _result_T_2170 = _result_T_2168 + _result_T_586;
  wire [63:0] _result_T_2172 = _result_T_2170 + _result_T_587;
  wire [63:0] _result_T_2174 = _result_T_2172 + _result_T_588;
  wire [63:0] _result_T_2176 = _result_T_2174 + _result_T_589;
  wire [63:0] _result_T_2178 = _result_T_2176 + _result_T_590;
  wire [63:0] _result_T_2180 = _result_T_2178 + _result_T_591;
  wire [63:0] _result_T_2182 = _result_T_2180 + _result_T_592;
  wire [63:0] _result_T_2184 = _result_T_2182 + _result_T_593;
  wire [63:0] _result_T_2186 = _result_T_2184 + _result_T_594;
  wire [63:0] _result_T_2188 = _result_T_2186 + _result_T_595;
  wire [63:0] _result_T_2190 = _result_T_2188 + _result_T_596;
  wire [63:0] _result_T_2192 = _result_T_2190 + _result_T_597;
  wire [63:0] _result_T_2194 = _result_T_2192 + _result_T_598;
  wire [63:0] _result_T_2196 = _result_T_2194 + _result_T_599;
  wire [63:0] _result_T_2198 = _result_T_2196 + _result_T_600;
  wire [63:0] _result_T_2200 = _result_T_2198 + _result_T_601;
  wire [63:0] _result_T_2202 = _result_T_2200 + _result_T_602;
  wire [63:0] _result_T_2204 = _result_T_2202 + _result_T_603;
  wire [63:0] _result_T_2206 = _result_T_2204 + _result_T_604;
  wire [63:0] _result_T_2208 = _result_T_2206 + _result_T_605;
  wire [63:0] _result_T_2210 = _result_T_2208 + _result_T_606;
  wire [63:0] _result_T_2212 = _result_T_2210 + _result_T_607;
  wire [63:0] _result_T_2214 = _result_T_2212 + _result_T_608;
  wire [63:0] _result_T_2216 = _result_T_2214 + _result_T_609;
  wire [63:0] _result_T_2218 = _result_T_2216 + _result_T_610;
  wire [63:0] _result_T_2220 = _result_T_2218 + _result_T_611;
  wire [63:0] _result_T_2222 = _result_T_2220 + _result_T_612;
  wire [63:0] _result_T_2224 = _result_T_2222 + _result_T_613;
  wire [63:0] _result_T_2226 = _result_T_2224 + _result_T_614;
  wire [63:0] _result_T_2228 = _result_T_2226 + _result_T_615;
  wire [63:0] _result_T_2230 = _result_T_2228 + _result_T_616;
  wire [63:0] _result_T_2232 = _result_T_2230 + _result_T_617;
  wire [63:0] _result_T_2234 = _result_T_2232 + _result_T_618;
  wire [63:0] _result_T_2236 = _result_T_2234 + _result_T_619;
  wire [63:0] _result_T_2238 = _result_T_2236 + _result_T_620;
  wire [63:0] _result_T_2240 = _result_T_2238 + _result_T_621;
  wire [63:0] _result_T_2242 = _result_T_2240 + _result_T_622;
  wire [63:0] _result_T_2244 = _result_T_2242 + _result_T_623;
  wire [63:0] _result_T_2246 = _result_T_2244 + _result_T_624;
  wire [63:0] _result_T_2248 = _result_T_2246 + _result_T_625;
  wire [63:0] _result_T_2250 = _result_T_2248 + _result_T_626;
  wire [63:0] _result_T_2252 = _result_T_2250 + _result_T_627;
  wire [63:0] _result_T_2254 = _result_T_2252 + _result_T_628;
  wire [63:0] _result_T_2256 = _result_T_2254 + _result_T_629;
  wire [63:0] _result_T_2258 = _result_T_2256 + _result_T_630;
  wire [63:0] _result_T_2260 = _result_T_2258 + _result_T_631;
  wire [63:0] _result_T_2262 = _result_T_2260 + _result_T_632;
  wire [63:0] _result_T_2264 = _result_T_2262 + _result_T_633;
  wire [63:0] _result_T_2266 = _result_T_2264 + _result_T_634;
  wire [63:0] _result_T_2268 = _result_T_2266 + _result_T_635;
  wire [63:0] _result_T_2270 = _result_T_2268 + _result_T_636;
  wire [63:0] _result_T_2272 = _result_T_2270 + _result_T_637;
  wire [63:0] _result_T_2274 = _result_T_2272 + _result_T_638;
  wire [63:0] _result_T_2276 = _result_T_2274 + _result_T_639;
  wire [63:0] _result_T_2278 = _result_T_2276 + _result_T_640;
  wire [63:0] _result_T_2280 = _result_T_2278 + _result_T_641;
  wire [63:0] _result_T_2282 = _result_T_2280 + _result_T_642;
  wire [63:0] _result_T_2284 = _result_T_2282 + _result_T_643;
  wire [63:0] _result_T_2286 = _result_T_2284 + _result_T_644;
  wire [63:0] _result_T_2288 = _result_T_2286 + _result_T_645;
  wire [63:0] _result_T_2290 = _result_T_2288 + _result_T_646;
  wire [63:0] _result_T_2292 = _result_T_2290 + _result_T_647;
  wire [63:0] _result_T_2294 = _result_T_2292 + _result_T_648;
  wire [63:0] _result_T_2296 = _result_T_2294 + _result_T_649;
  wire [63:0] _result_T_2298 = _result_T_2296 + _result_T_650;
  wire [63:0] _result_T_2300 = _result_T_2298 + _result_T_651;
  wire [63:0] _result_T_2302 = _result_T_2300 + _result_T_652;
  wire [63:0] _result_T_2304 = _result_T_2302 + _result_T_653;
  wire [63:0] _result_T_2306 = _result_T_2304 + _result_T_654;
  wire [63:0] _result_T_2308 = _result_T_2306 + _result_T_655;
  wire [63:0] _result_T_2310 = _result_T_2308 + _result_T_656;
  wire [63:0] _result_T_2312 = _result_T_2310 + _result_T_657;
  wire [63:0] _result_T_2314 = _result_T_2312 + _result_T_658;
  wire [63:0] _result_T_2316 = _result_T_2314 + _result_T_659;
  wire [63:0] _result_T_2318 = _result_T_2316 + _result_T_660;
  wire [63:0] _result_T_2320 = _result_T_2318 + _result_T_661;
  wire [63:0] _result_T_2322 = _result_T_2320 + _result_T_662;
  wire [63:0] _result_T_2324 = _result_T_2322 + _result_T_663;
  wire [63:0] _result_T_2326 = _result_T_2324 + _result_T_664;
  wire [63:0] _result_T_2328 = _result_T_2326 + _result_T_665;
  wire [63:0] _result_T_2330 = _result_T_2328 + _result_T_666;
  wire [63:0] _result_T_2332 = _result_T_2330 + _result_T_667;
  wire [63:0] _result_T_2334 = _result_T_2332 + _result_T_668;
  wire [63:0] _result_T_2336 = _result_T_2334 + _result_T_669;
  wire [63:0] _result_T_2338 = _result_T_2336 + _result_T_670;
  wire [63:0] _result_T_2340 = _result_T_2338 + _result_T_671;
  wire [63:0] _result_T_2342 = _result_T_2340 + _result_T_672;
  wire [63:0] _result_T_2344 = _result_T_2342 + _result_T_673;
  wire [63:0] _result_T_2346 = _result_T_2344 + _result_T_674;
  wire [63:0] _result_T_2348 = _result_T_2346 + _result_T_675;
  wire [63:0] _result_T_2350 = _result_T_2348 + _result_T_676;
  wire [63:0] _result_T_2352 = _result_T_2350 + _result_T_677;
  wire [63:0] _result_T_2354 = _result_T_2352 + _result_T_678;
  wire [63:0] _result_T_2356 = _result_T_2354 + _result_T_679;
  wire [63:0] _result_T_2358 = _result_T_2356 + _result_T_680;
  wire [63:0] _result_T_2360 = _result_T_2358 + _result_T_681;
  wire [63:0] _result_T_2362 = _result_T_2360 + _result_T_682;
  wire [63:0] _result_T_2364 = _result_T_2362 + _result_T_683;
  wire [63:0] _result_T_2366 = _result_T_2364 + _result_T_684;
  wire [63:0] _result_T_2368 = _result_T_2366 + _result_T_685;
  wire [63:0] _result_T_2370 = _result_T_2368 + _result_T_686;
  wire [63:0] _result_T_2372 = _result_T_2370 + _result_T_687;
  wire [63:0] _result_T_2374 = _result_T_2372 + _result_T_688;
  wire [63:0] _result_T_2376 = _result_T_2374 + _result_T_689;
  wire [63:0] _result_T_2378 = _result_T_2376 + _result_T_690;
  wire [63:0] _result_T_2380 = _result_T_2378 + _result_T_691;
  wire [63:0] _result_T_2382 = _result_T_2380 + _result_T_692;
  wire [63:0] _result_T_2384 = _result_T_2382 + _result_T_693;
  wire [63:0] _result_T_2386 = _result_T_2384 + _result_T_694;
  wire [63:0] _result_T_2388 = _result_T_2386 + _result_T_695;
  wire [63:0] _result_T_2390 = _result_T_2388 + _result_T_696;
  wire [63:0] _result_T_2392 = _result_T_2390 + _result_T_697;
  wire [63:0] _result_T_2394 = _result_T_2392 + _result_T_698;
  wire [63:0] _result_T_2396 = _result_T_2394 + _result_T_699;
  wire [63:0] _result_T_2398 = _result_T_2396 + _result_T_700;
  wire [63:0] _result_T_2400 = _result_T_2398 + _result_T_701;
  wire [63:0] _result_T_2402 = _result_T_2400 + _result_T_702;
  wire [63:0] _result_T_2404 = _result_T_2402 + _result_T_703;
  wire [63:0] _result_T_2406 = _result_T_2404 + _result_T_704;
  wire [63:0] _result_T_2408 = _result_T_2406 + _result_T_705;
  wire [63:0] _result_T_2410 = _result_T_2408 + _result_T_706;
  wire [63:0] _result_T_2412 = _result_T_2410 + _result_T_707;
  wire [63:0] _result_T_2414 = _result_T_2412 + _result_T_708;
  wire [63:0] _result_T_2416 = _result_T_2414 + _result_T_709;
  wire [63:0] _result_T_2418 = _result_T_2416 + _result_T_710;
  wire [63:0] _result_T_2420 = _result_T_2418 + _result_T_711;
  wire [63:0] _result_T_2422 = _result_T_2420 + _result_T_712;
  wire [63:0] _result_T_2424 = _result_T_2422 + _result_T_713;
  wire [63:0] _result_T_2426 = _result_T_2424 + _result_T_714;
  wire [63:0] _result_T_2428 = _result_T_2426 + _result_T_715;
  wire [63:0] _result_T_2430 = _result_T_2428 + _result_T_716;
  wire [63:0] _result_T_2432 = _result_T_2430 + _result_T_717;
  wire [63:0] _result_T_2434 = _result_T_2432 + _result_T_718;
  wire [63:0] _result_T_2436 = _result_T_2434 + _result_T_719;
  wire [63:0] _result_T_2438 = _result_T_2436 + _result_T_720;
  wire [63:0] _result_T_2440 = _result_T_2438 + _result_T_721;
  wire [63:0] _result_T_2442 = _result_T_2440 + _result_T_722;
  wire [63:0] _result_T_2444 = _result_T_2442 + _result_T_723;
  wire [63:0] _result_T_2446 = _result_T_2444 + _result_T_724;
  wire [63:0] _result_T_2448 = _result_T_2446 + _result_T_725;
  wire [63:0] _result_T_2450 = _result_T_2448 + _result_T_726;
  wire [63:0] _result_T_2452 = _result_T_2450 + _result_T_727;
  wire [63:0] _result_T_2454 = _result_T_2452 + _result_T_728;
  wire [63:0] _result_T_2456 = _result_T_2454 + _result_T_729;
  wire [63:0] _result_T_2458 = _result_T_2456 + _result_T_730;
  wire [63:0] _result_T_2460 = _result_T_2458 + _result_T_731;
  wire [63:0] _result_T_2462 = _result_T_2460 + _result_T_732;
  wire [63:0] _result_T_2464 = _result_T_2462 + _result_T_733;
  wire [63:0] _result_T_2466 = _result_T_2464 + _result_T_734;
  wire [63:0] _result_T_2468 = _result_T_2466 + _result_T_735;
  wire [63:0] _result_T_2470 = _result_T_2468 + _result_T_736;
  wire [63:0] _result_T_2472 = _result_T_2470 + _result_T_737;
  wire [63:0] _result_T_2474 = _result_T_2472 + _result_T_738;
  wire [63:0] _result_T_2476 = _result_T_2474 + _result_T_739;
  wire [63:0] _result_T_2478 = _result_T_2476 + _result_T_740;
  wire [63:0] _result_T_2480 = _result_T_2478 + _result_T_741;
  wire [63:0] _result_T_2482 = _result_T_2480 + _result_T_742;
  wire [63:0] _result_T_2484 = _result_T_2482 + _result_T_743;
  wire [63:0] _result_T_2486 = _result_T_2484 + _result_T_744;
  wire [63:0] _result_T_2488 = _result_T_2486 + _result_T_745;
  wire [63:0] _result_T_2490 = _result_T_2488 + _result_T_746;
  wire [63:0] _result_T_2492 = _result_T_2490 + _result_T_747;
  wire [63:0] _result_T_2494 = _result_T_2492 + _result_T_748;
  wire [63:0] _result_T_2496 = _result_T_2494 + _result_T_749;
  wire [63:0] _result_T_2498 = _result_T_2496 + _result_T_750;
  wire [63:0] _result_T_2500 = _result_T_2498 + _result_T_751;
  wire [63:0] _result_T_2502 = _result_T_2500 + _result_T_752;
  wire [63:0] _result_T_2504 = _result_T_2502 + _result_T_753;
  wire [63:0] _result_T_2506 = _result_T_2504 + _result_T_754;
  wire [63:0] _result_T_2508 = _result_T_2506 + _result_T_755;
  wire [63:0] _result_T_2510 = _result_T_2508 + _result_T_756;
  wire [63:0] _result_T_2512 = _result_T_2510 + _result_T_757;
  wire [63:0] _result_T_2514 = _result_T_2512 + _result_T_758;
  wire [63:0] _result_T_2516 = _result_T_2514 + _result_T_759;
  wire [63:0] _result_T_2518 = _result_T_2516 + _result_T_760;
  wire [63:0] _result_T_2520 = _result_T_2518 + _result_T_761;
  wire [63:0] _result_T_2522 = _result_T_2520 + _result_T_762;
  wire [63:0] _result_T_2524 = _result_T_2522 + _result_T_763;
  wire [63:0] _result_T_2526 = _result_T_2524 + _result_T_764;
  wire [63:0] _result_T_2528 = _result_T_2526 + _result_T_765;
  wire [63:0] _result_T_2530 = _result_T_2528 + _result_T_766;
  wire [63:0] _result_T_2532 = _result_T_2530 + _result_T_767;
  wire [63:0] _result_T_2534 = _result_T_2532 + _result_T_768;
  wire [63:0] _result_T_2536 = _result_T_2534 + _result_T_769;
  wire [63:0] _result_T_2538 = _result_T_2536 + _result_T_770;
  wire [63:0] _result_T_2540 = _result_T_2538 + _result_T_771;
  wire [63:0] _result_T_2542 = _result_T_2540 + _result_T_772;
  wire [63:0] _result_T_2544 = _result_T_2542 + _result_T_773;
  wire [63:0] _result_T_2546 = _result_T_2544 + _result_T_774;
  wire [63:0] _result_T_2548 = _result_T_2546 + _result_T_775;
  wire [63:0] _result_T_2550 = _result_T_2548 + _result_T_776;
  wire [63:0] _result_T_2552 = _result_T_2550 + _result_T_777;
  wire [63:0] _result_T_2554 = _result_T_2552 + _result_T_778;
  wire [63:0] _result_T_2556 = _result_T_2554 + _result_T_779;
  wire [63:0] _result_T_2558 = _result_T_2556 + _result_T_780;
  wire [63:0] _result_T_2560 = _result_T_2558 + _result_T_781;
  wire [63:0] _result_T_2562 = _result_T_2560 + _result_T_782;
  wire [63:0] _result_T_2564 = _result_T_2562 + _result_T_783;
  wire [63:0] _result_T_2566 = _result_T_2564 + _result_T_784;
  wire [63:0] _result_T_2568 = _result_T_2566 + _result_T_785;
  wire [63:0] _result_T_2570 = _result_T_2568 + _result_T_786;
  wire [63:0] _result_T_2572 = _result_T_2570 + _result_T_787;
  wire [63:0] _result_T_2574 = _result_T_2572 + _result_T_788;
  wire [63:0] _result_T_2576 = _result_T_2574 + _result_T_789;
  wire [63:0] _result_T_2578 = _result_T_2576 + _result_T_790;
  wire [63:0] _result_T_2580 = _result_T_2578 + _result_T_791;
  wire [63:0] _result_T_2582 = _result_T_2580 + _result_T_792;
  wire [63:0] _result_T_2584 = _result_T_2582 + _result_T_793;
  wire [63:0] _result_T_2586 = _result_T_2584 + _result_T_794;
  wire [63:0] _result_T_2588 = _result_T_2586 + _result_T_795;
  wire [63:0] _result_T_2590 = _result_T_2588 + _result_T_796;
  wire [63:0] _result_T_2592 = _result_T_2590 + _result_T_797;
  wire [63:0] _result_T_2594 = _result_T_2592 + _result_T_798;
  wire [63:0] _result_T_2596 = _result_T_2594 + _result_T_799;
  wire [63:0] _result_T_2598 = _result_T_2596 + _result_T_800;
  wire [63:0] _result_T_2600 = _result_T_2598 + _result_T_801;
  wire [63:0] _result_T_2602 = _result_T_2600 + _result_T_802;
  wire [63:0] _result_T_2604 = _result_T_2602 + _result_T_803;
  wire [63:0] _result_T_2606 = _result_T_2604 + _result_T_804;
  wire [63:0] _result_T_2608 = _result_T_2606 + _result_T_805;
  wire [63:0] _result_T_2610 = _result_T_2608 + _result_T_806;
  wire [63:0] _result_T_2612 = _result_T_2610 + _result_T_807;
  wire [63:0] _result_T_2614 = _result_T_2612 + _result_T_808;
  wire [63:0] _result_T_2616 = _result_T_2614 + _result_T_809;
  wire [63:0] _result_T_2618 = _result_T_2616 + _result_T_810;
  wire [63:0] _result_T_2620 = _result_T_2618 + _result_T_811;
  wire [63:0] _result_T_2622 = _result_T_2620 + _result_T_812;
  wire [63:0] _result_T_2624 = _result_T_2622 + _result_T_813;
  wire [63:0] _result_T_2626 = _result_T_2624 + _result_T_814;
  wire [63:0] _result_T_2628 = _result_T_2626 + _result_T_815;
  wire [63:0] _result_T_2630 = _result_T_2628 + _result_T_816;
  wire [63:0] _result_T_2632 = _result_T_2630 + _result_T_817;
  wire [63:0] _result_T_2634 = _result_T_2632 + _result_T_818;
  wire [63:0] _result_T_2636 = _result_T_2634 + _result_T_819;
  wire [63:0] _result_T_2638 = _result_T_2636 + _result_T_820;
  wire [63:0] _result_T_2640 = _result_T_2638 + _result_T_821;
  wire [63:0] _result_T_2642 = _result_T_2640 + _result_T_822;
  wire [63:0] _result_T_2644 = _result_T_2642 + _result_T_823;
  wire [63:0] _result_T_2646 = _result_T_2644 + _result_T_824;
  wire [63:0] _result_T_2648 = _result_T_2646 + _result_T_825;
  wire [63:0] _result_T_2650 = _result_T_2648 + _result_T_826;
  wire [63:0] _result_T_2652 = _result_T_2650 + _result_T_827;
  wire [63:0] _result_T_2654 = _result_T_2652 + _result_T_828;
  wire [63:0] _result_T_2656 = _result_T_2654 + _result_T_829;
  wire [63:0] _result_T_2658 = _result_T_2656 + _result_T_830;
  wire [63:0] _result_T_2660 = _result_T_2658 + _result_T_831;
  wire [63:0] _result_T_2662 = _result_T_2660 + _result_T_832;
  wire [63:0] _result_T_2664 = _result_T_2662 + _result_T_833;
  wire [63:0] _result_T_2666 = _result_T_2664 + _result_T_834;
  wire [63:0] _result_T_2668 = _result_T_2666 + _result_T_835;
  wire [63:0] _result_T_2670 = _result_T_2668 + _result_T_836;
  wire [63:0] _result_T_2672 = _result_T_2670 + _result_T_837;
  wire [63:0] _result_T_2674 = _result_T_2672 + _result_T_838;
  wire [63:0] _result_T_2676 = _result_T_2674 + _result_T_839;
  wire [63:0] _result_T_2678 = _result_T_2676 + _result_T_840;
  wire [63:0] _result_T_2680 = _result_T_2678 + _result_T_841;
  wire [63:0] _result_T_2682 = _result_T_2680 + _result_T_842;
  wire [63:0] _result_T_2684 = _result_T_2682 + _result_T_843;
  wire [63:0] _result_T_2686 = _result_T_2684 + _result_T_844;
  wire [63:0] _result_T_2688 = _result_T_2686 + _result_T_845;
  wire [63:0] _result_T_2690 = _result_T_2688 + _result_T_846;
  wire [63:0] _result_T_2692 = _result_T_2690 + _result_T_847;
  wire [63:0] _result_T_2694 = _result_T_2692 + _result_T_848;
  wire [63:0] _result_T_2696 = _result_T_2694 + _result_T_849;
  wire [63:0] _result_T_2698 = _result_T_2696 + _result_T_850;
  wire [63:0] _result_T_2700 = _result_T_2698 + _result_T_851;
  wire [63:0] _result_T_2702 = _result_T_2700 + _result_T_852;
  wire [63:0] _result_T_2704 = _result_T_2702 + _result_T_853;
  wire [63:0] _result_T_2706 = _result_T_2704 + _result_T_854;
  wire [63:0] _result_T_2708 = _result_T_2706 + _result_T_855;
  wire [63:0] _result_T_2710 = _result_T_2708 + _result_T_856;
  wire [63:0] _result_T_2712 = _result_T_2710 + _result_T_857;
  wire [63:0] _result_T_2714 = _result_T_2712 + _result_T_858;
  wire [63:0] _result_T_2716 = _result_T_2714 + _result_T_859;
  wire [63:0] _result_T_2718 = _result_T_2716 + _result_T_860;
  wire [63:0] _result_T_2720 = _result_T_2718 + _result_T_861;
  wire [63:0] _result_T_2722 = _result_T_2720 + _result_T_862;
  wire [63:0] _result_T_2724 = _result_T_2722 + _result_T_863;
  wire [63:0] _result_T_2726 = _result_T_2724 + _result_T_864;
  wire [63:0] _result_T_2728 = _result_T_2726 + _result_T_865;
  wire [63:0] _result_T_2730 = _result_T_2728 + _result_T_866;
  wire [63:0] _result_T_2732 = _result_T_2730 + _result_T_867;
  wire [63:0] _result_T_2734 = _result_T_2732 + _result_T_868;
  wire [63:0] _result_T_2736 = _result_T_2734 + _result_T_869;
  wire [63:0] _result_T_2738 = _result_T_2736 + _result_T_870;
  wire [63:0] _result_T_2740 = _result_T_2738 + _result_T_871;
  wire [63:0] _result_T_2742 = _result_T_2740 + _result_T_872;
  wire [63:0] _result_T_2744 = _result_T_2742 + _result_T_873;
  wire [63:0] _result_T_2746 = _result_T_2744 + _result_T_874;
  wire [63:0] _result_T_2748 = _result_T_2746 + _result_T_875;
  wire [63:0] _result_T_2750 = _result_T_2748 + _result_T_876;
  wire [63:0] _result_T_2752 = _result_T_2750 + _result_T_877;
  wire [63:0] _result_T_2754 = _result_T_2752 + _result_T_878;
  wire [63:0] _result_T_2756 = _result_T_2754 + _result_T_879;
  wire [63:0] _result_T_2758 = _result_T_2756 + _result_T_880;
  wire [63:0] _result_T_2760 = _result_T_2758 + _result_T_881;
  wire [63:0] _result_T_2762 = _result_T_2760 + _result_T_882;
  wire [63:0] _result_T_2764 = _result_T_2762 + _result_T_883;
  wire [63:0] _result_T_2766 = _result_T_2764 + _result_T_884;
  wire [63:0] _result_T_2768 = _result_T_2766 + _result_T_885;
  wire [63:0] _result_T_2770 = _result_T_2768 + _result_T_886;
  wire [63:0] _result_T_2772 = _result_T_2770 + _result_T_887;
  wire [63:0] _result_T_2774 = _result_T_2772 + _result_T_888;
  wire [63:0] _result_T_2776 = _result_T_2774 + _result_T_889;
  wire [63:0] _result_T_2778 = _result_T_2776 + _result_T_890;
  wire [63:0] _result_T_2780 = _result_T_2778 + _result_T_891;
  wire [63:0] _result_T_2782 = _result_T_2780 + _result_T_892;
  wire [63:0] _result_T_2784 = _result_T_2782 + _result_T_893;
  wire [63:0] _result_T_2786 = _result_T_2784 + _result_T_894;
  wire [63:0] _result_T_2788 = _result_T_2786 + _result_T_895;
  wire [63:0] _result_T_2790 = _result_T_2788 + _result_T_896;
  wire [63:0] _result_T_2792 = _result_T_2790 + _result_T_897;
  wire [63:0] _result_T_2794 = _result_T_2792 + _result_T_898;
  wire [63:0] _result_T_2796 = _result_T_2794 + _result_T_899;
  wire [63:0] _result_T_2798 = _result_T_2796 + _result_T_900;
  wire [63:0] _result_T_2800 = _result_T_2798 + _result_T_901;
  wire [63:0] _result_T_2802 = _result_T_2800 + _result_T_902;
  wire [63:0] _result_T_2804 = _result_T_2802 + _result_T_903;
  wire [63:0] _result_T_2806 = _result_T_2804 + _result_T_904;
  wire [63:0] _result_T_2808 = _result_T_2806 + _result_T_905;
  wire [63:0] _result_T_2810 = _result_T_2808 + _result_T_906;
  wire [63:0] _result_T_2812 = _result_T_2810 + _result_T_907;
  wire [63:0] _result_T_2814 = _result_T_2812 + _result_T_908;
  wire [63:0] _result_T_2816 = _result_T_2814 + _result_T_909;
  wire [63:0] _result_T_2818 = _result_T_2816 + _result_T_910;
  wire [63:0] _result_T_2820 = _result_T_2818 + _result_T_911;
  wire [63:0] _result_T_2822 = _result_T_2820 + _result_T_912;
  wire [63:0] _result_T_2824 = _result_T_2822 + _result_T_913;
  wire [63:0] _result_T_2826 = _result_T_2824 + _result_T_914;
  wire [63:0] _result_T_2828 = _result_T_2826 + _result_T_915;
  wire [63:0] _result_T_2830 = _result_T_2828 + _result_T_916;
  wire [63:0] _result_T_2832 = _result_T_2830 + _result_T_917;
  wire [63:0] _result_T_2834 = _result_T_2832 + _result_T_918;
  wire [63:0] _result_T_2836 = _result_T_2834 + _result_T_919;
  wire [63:0] _result_T_2838 = _result_T_2836 + _result_T_920;
  wire [63:0] _result_T_2840 = _result_T_2838 + _result_T_921;
  wire [63:0] _result_T_2842 = _result_T_2840 + _result_T_922;
  wire [63:0] _result_T_2844 = _result_T_2842 + _result_T_923;
  wire [63:0] _result_T_2846 = _result_T_2844 + _result_T_924;
  wire [63:0] _result_T_2848 = _result_T_2846 + _result_T_925;
  wire [63:0] _result_T_2850 = _result_T_2848 + _result_T_926;
  wire [63:0] _result_T_2852 = _result_T_2850 + _result_T_927;
  wire [63:0] _result_T_2854 = _result_T_2852 + _result_T_928;
  wire [63:0] _result_T_2856 = _result_T_2854 + _result_T_929;
  wire [63:0] _result_T_2858 = _result_T_2856 + _result_T_930;
  wire [63:0] _result_T_2860 = _result_T_2858 + _result_T_931;
  wire [63:0] _result_T_2862 = _result_T_2860 + _result_T_932;
  wire [63:0] _result_T_2864 = _result_T_2862 + _result_T_933;
  wire [63:0] _result_T_2866 = _result_T_2864 + _result_T_934;
  wire [63:0] _result_T_2868 = _result_T_2866 + _result_T_935;
  wire [63:0] _result_T_2870 = _result_T_2868 + _result_T_936;
  wire [63:0] _result_T_2872 = _result_T_2870 + _result_T_937;
  wire [63:0] _result_T_2874 = _result_T_2872 + _result_T_938;
  wire [63:0] _result_T_2876 = _result_T_2874 + _result_T_939;
  wire [63:0] _result_T_2878 = _result_T_2876 + _result_T_940;
  wire [63:0] _result_T_2880 = _result_T_2878 + _result_T_941;
  wire [63:0] _result_T_2882 = _result_T_2880 + _result_T_942;
  wire [63:0] _result_T_2884 = _result_T_2882 + _result_T_943;
  wire [63:0] _result_T_2886 = _result_T_2884 + _result_T_944;
  wire [63:0] _result_T_2888 = _result_T_2886 + _result_T_945;
  wire [63:0] _result_T_2890 = _result_T_2888 + _result_T_946;
  wire [63:0] _result_T_2892 = _result_T_2890 + _result_T_947;
  wire [63:0] _result_T_2894 = _result_T_2892 + _result_T_948;
  wire [63:0] _result_T_2896 = _result_T_2894 + _result_T_949;
  wire [63:0] _result_T_2898 = _result_T_2896 + _result_T_950;
  wire [63:0] _result_T_2900 = _result_T_2898 + _result_T_951;
  wire [63:0] _result_T_2902 = _result_T_2900 + _result_T_952;
  wire [63:0] _result_T_2904 = _result_T_2902 + _result_T_953;
  wire [63:0] _result_T_2906 = _result_T_2904 + _result_T_954;
  wire [63:0] _result_T_2908 = _result_T_2906 + _result_T_955;
  wire [63:0] _result_T_2910 = _result_T_2908 + _result_T_956;
  wire [63:0] _result_T_2912 = _result_T_2910 + _result_T_957;
  wire [63:0] _result_T_2914 = _result_T_2912 + _result_T_958;
  wire [63:0] _result_T_2916 = _result_T_2914 + _result_T_959;
  wire [63:0] _result_T_2918 = _result_T_2916 + _result_T_960;
  wire [63:0] _result_T_2920 = _result_T_2918 + _result_T_961;
  wire [63:0] _result_T_2922 = _result_T_2920 + _result_T_962;
  wire [63:0] _result_T_2924 = _result_T_2922 + _result_T_963;
  wire [63:0] _result_T_2926 = _result_T_2924 + _result_T_964;
  wire [63:0] _result_T_2928 = _result_T_2926 + _result_T_965;
  wire [63:0] _result_T_2930 = _result_T_2928 + _result_T_966;
  wire [63:0] _result_T_2932 = _result_T_2930 + _result_T_967;
  wire [63:0] _result_T_2934 = _result_T_2932 + _result_T_968;
  wire [63:0] _result_T_2936 = _result_T_2934 + _result_T_969;
  wire [63:0] _result_T_2938 = _result_T_2936 + _result_T_970;
  wire [63:0] _result_T_2940 = _result_T_2938 + _result_T_971;
  wire [63:0] _result_T_2942 = _result_T_2940 + _result_T_972;
  wire [63:0] _result_T_2944 = _result_T_2942 + _result_T_973;
  wire [63:0] _result_T_2946 = _result_T_2944 + _result_T_974;
  wire [63:0] _result_T_2948 = _result_T_2946 + _result_T_975;
  wire [63:0] _result_T_2950 = _result_T_2948 + _result_T_976;
  wire [63:0] _result_T_2952 = _result_T_2950 + _result_T_977;
  wire [63:0] _result_T_2954 = _result_T_2952 + _result_T_978;
  wire [63:0] _result_T_2956 = _result_T_2954 + _result_T_979;
  wire [63:0] _result_T_2958 = _result_T_2956 + _result_T_980;
  wire [63:0] _result_T_2960 = _result_T_2958 + _result_T_981;
  wire [63:0] _result_T_2962 = _result_T_2960 + _result_T_982;
  wire [63:0] _result_T_2964 = _result_T_2962 + _result_T_983;
  wire [63:0] _result_T_2966 = _result_T_2964 + _result_T_984;
  wire [63:0] _result_T_2968 = _result_T_2966 + _result_T_985;
  wire [63:0] _result_T_2970 = _result_T_2968 + _result_T_986;
  wire [63:0] _result_T_2972 = _result_T_2970 + _result_T_987;
  wire [63:0] _result_T_2974 = _result_T_2972 + _result_T_988;
  wire [63:0] _result_T_2976 = _result_T_2974 + _result_T_989;
  wire [63:0] _result_T_2978 = _result_T_2976 + _result_T_990;
  wire [63:0] _result_T_2980 = _result_T_2978 + _result_T_991;
  wire [63:0] _result_T_2982 = _result_T_2980 + _result_T_992;
  wire [63:0] _result_T_2984 = _result_T_2982 + _result_T_993;
  wire [63:0] _result_T_2986 = _result_T_2984 + _result_T_994;
  wire [63:0] _result_T_2988 = _result_T_2986 + _result_T_995;
  wire [63:0] _result_T_2990 = _result_T_2988 + _result_T_996;
  wire [63:0] _result_T_2992 = _result_T_2990 + _result_T_997;
  wire [63:0] _result_T_2994 = _result_T_2992 + _result_T_998;
  wire [63:0] _result_T_2996 = _result_T_2994 + _result_T_999;
  wire [63:0] _result_T_2998 = _result_T_2996 + _result_T_1000;
  wire [63:0] _GEN_2000 = insn[6:0] == 7'h3b ? _result_T_2998 : result;
  assign rd = result[31:0];
  always @(posedge clock) begin
    if (reset) begin
      coeffs_0 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h0 == rs2[9:0]) begin
          coeffs_0 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_1 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1 == rs2[9:0]) begin
          coeffs_1 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_2 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2 == rs2[9:0]) begin
          coeffs_2 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_3 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3 == rs2[9:0]) begin
          coeffs_3 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_4 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h4 == rs2[9:0]) begin
          coeffs_4 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_5 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h5 == rs2[9:0]) begin
          coeffs_5 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_6 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h6 == rs2[9:0]) begin
          coeffs_6 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_7 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h7 == rs2[9:0]) begin
          coeffs_7 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_8 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h8 == rs2[9:0]) begin
          coeffs_8 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_9 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h9 == rs2[9:0]) begin
          coeffs_9 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_10 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha == rs2[9:0]) begin
          coeffs_10 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_11 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb == rs2[9:0]) begin
          coeffs_11 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_12 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc == rs2[9:0]) begin
          coeffs_12 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_13 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd == rs2[9:0]) begin
          coeffs_13 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_14 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he == rs2[9:0]) begin
          coeffs_14 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_15 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf == rs2[9:0]) begin
          coeffs_15 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_16 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h10 == rs2[9:0]) begin
          coeffs_16 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_17 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h11 == rs2[9:0]) begin
          coeffs_17 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_18 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h12 == rs2[9:0]) begin
          coeffs_18 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_19 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h13 == rs2[9:0]) begin
          coeffs_19 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_20 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h14 == rs2[9:0]) begin
          coeffs_20 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_21 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h15 == rs2[9:0]) begin
          coeffs_21 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_22 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h16 == rs2[9:0]) begin
          coeffs_22 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_23 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h17 == rs2[9:0]) begin
          coeffs_23 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_24 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h18 == rs2[9:0]) begin
          coeffs_24 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_25 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h19 == rs2[9:0]) begin
          coeffs_25 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_26 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a == rs2[9:0]) begin
          coeffs_26 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_27 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b == rs2[9:0]) begin
          coeffs_27 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_28 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c == rs2[9:0]) begin
          coeffs_28 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_29 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d == rs2[9:0]) begin
          coeffs_29 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_30 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e == rs2[9:0]) begin
          coeffs_30 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_31 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f == rs2[9:0]) begin
          coeffs_31 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_32 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h20 == rs2[9:0]) begin
          coeffs_32 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_33 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h21 == rs2[9:0]) begin
          coeffs_33 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_34 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h22 == rs2[9:0]) begin
          coeffs_34 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_35 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h23 == rs2[9:0]) begin
          coeffs_35 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_36 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h24 == rs2[9:0]) begin
          coeffs_36 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_37 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h25 == rs2[9:0]) begin
          coeffs_37 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_38 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h26 == rs2[9:0]) begin
          coeffs_38 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_39 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h27 == rs2[9:0]) begin
          coeffs_39 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_40 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h28 == rs2[9:0]) begin
          coeffs_40 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_41 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h29 == rs2[9:0]) begin
          coeffs_41 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_42 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a == rs2[9:0]) begin
          coeffs_42 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_43 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b == rs2[9:0]) begin
          coeffs_43 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_44 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c == rs2[9:0]) begin
          coeffs_44 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_45 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d == rs2[9:0]) begin
          coeffs_45 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_46 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e == rs2[9:0]) begin
          coeffs_46 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_47 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f == rs2[9:0]) begin
          coeffs_47 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_48 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h30 == rs2[9:0]) begin
          coeffs_48 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_49 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h31 == rs2[9:0]) begin
          coeffs_49 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_50 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h32 == rs2[9:0]) begin
          coeffs_50 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_51 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h33 == rs2[9:0]) begin
          coeffs_51 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_52 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h34 == rs2[9:0]) begin
          coeffs_52 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_53 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h35 == rs2[9:0]) begin
          coeffs_53 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_54 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h36 == rs2[9:0]) begin
          coeffs_54 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_55 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h37 == rs2[9:0]) begin
          coeffs_55 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_56 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h38 == rs2[9:0]) begin
          coeffs_56 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_57 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h39 == rs2[9:0]) begin
          coeffs_57 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_58 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a == rs2[9:0]) begin
          coeffs_58 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_59 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b == rs2[9:0]) begin
          coeffs_59 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_60 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c == rs2[9:0]) begin
          coeffs_60 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_61 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d == rs2[9:0]) begin
          coeffs_61 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_62 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3e == rs2[9:0]) begin
          coeffs_62 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_63 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3f == rs2[9:0]) begin
          coeffs_63 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_64 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h40 == rs2[9:0]) begin
          coeffs_64 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_65 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h41 == rs2[9:0]) begin
          coeffs_65 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_66 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h42 == rs2[9:0]) begin
          coeffs_66 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_67 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h43 == rs2[9:0]) begin
          coeffs_67 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_68 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h44 == rs2[9:0]) begin
          coeffs_68 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_69 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h45 == rs2[9:0]) begin
          coeffs_69 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_70 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h46 == rs2[9:0]) begin
          coeffs_70 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_71 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h47 == rs2[9:0]) begin
          coeffs_71 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_72 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h48 == rs2[9:0]) begin
          coeffs_72 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_73 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h49 == rs2[9:0]) begin
          coeffs_73 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_74 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h4a == rs2[9:0]) begin
          coeffs_74 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_75 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h4b == rs2[9:0]) begin
          coeffs_75 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_76 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h4c == rs2[9:0]) begin
          coeffs_76 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_77 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h4d == rs2[9:0]) begin
          coeffs_77 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_78 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h4e == rs2[9:0]) begin
          coeffs_78 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_79 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h4f == rs2[9:0]) begin
          coeffs_79 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_80 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h50 == rs2[9:0]) begin
          coeffs_80 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_81 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h51 == rs2[9:0]) begin
          coeffs_81 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_82 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h52 == rs2[9:0]) begin
          coeffs_82 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_83 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h53 == rs2[9:0]) begin
          coeffs_83 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_84 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h54 == rs2[9:0]) begin
          coeffs_84 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_85 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h55 == rs2[9:0]) begin
          coeffs_85 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_86 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h56 == rs2[9:0]) begin
          coeffs_86 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_87 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h57 == rs2[9:0]) begin
          coeffs_87 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_88 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h58 == rs2[9:0]) begin
          coeffs_88 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_89 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h59 == rs2[9:0]) begin
          coeffs_89 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_90 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h5a == rs2[9:0]) begin
          coeffs_90 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_91 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h5b == rs2[9:0]) begin
          coeffs_91 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_92 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h5c == rs2[9:0]) begin
          coeffs_92 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_93 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h5d == rs2[9:0]) begin
          coeffs_93 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_94 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h5e == rs2[9:0]) begin
          coeffs_94 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_95 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h5f == rs2[9:0]) begin
          coeffs_95 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_96 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h60 == rs2[9:0]) begin
          coeffs_96 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_97 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h61 == rs2[9:0]) begin
          coeffs_97 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_98 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h62 == rs2[9:0]) begin
          coeffs_98 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_99 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h63 == rs2[9:0]) begin
          coeffs_99 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_100 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h64 == rs2[9:0]) begin
          coeffs_100 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_101 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h65 == rs2[9:0]) begin
          coeffs_101 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_102 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h66 == rs2[9:0]) begin
          coeffs_102 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_103 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h67 == rs2[9:0]) begin
          coeffs_103 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_104 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h68 == rs2[9:0]) begin
          coeffs_104 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_105 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h69 == rs2[9:0]) begin
          coeffs_105 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_106 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h6a == rs2[9:0]) begin
          coeffs_106 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_107 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h6b == rs2[9:0]) begin
          coeffs_107 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_108 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h6c == rs2[9:0]) begin
          coeffs_108 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_109 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h6d == rs2[9:0]) begin
          coeffs_109 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_110 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h6e == rs2[9:0]) begin
          coeffs_110 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_111 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h6f == rs2[9:0]) begin
          coeffs_111 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_112 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h70 == rs2[9:0]) begin
          coeffs_112 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_113 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h71 == rs2[9:0]) begin
          coeffs_113 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_114 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h72 == rs2[9:0]) begin
          coeffs_114 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_115 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h73 == rs2[9:0]) begin
          coeffs_115 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_116 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h74 == rs2[9:0]) begin
          coeffs_116 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_117 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h75 == rs2[9:0]) begin
          coeffs_117 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_118 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h76 == rs2[9:0]) begin
          coeffs_118 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_119 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h77 == rs2[9:0]) begin
          coeffs_119 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_120 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h78 == rs2[9:0]) begin
          coeffs_120 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_121 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h79 == rs2[9:0]) begin
          coeffs_121 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_122 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h7a == rs2[9:0]) begin
          coeffs_122 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_123 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h7b == rs2[9:0]) begin
          coeffs_123 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_124 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h7c == rs2[9:0]) begin
          coeffs_124 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_125 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h7d == rs2[9:0]) begin
          coeffs_125 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_126 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h7e == rs2[9:0]) begin
          coeffs_126 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_127 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h7f == rs2[9:0]) begin
          coeffs_127 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_128 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h80 == rs2[9:0]) begin
          coeffs_128 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_129 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h81 == rs2[9:0]) begin
          coeffs_129 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_130 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h82 == rs2[9:0]) begin
          coeffs_130 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_131 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h83 == rs2[9:0]) begin
          coeffs_131 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_132 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h84 == rs2[9:0]) begin
          coeffs_132 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_133 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h85 == rs2[9:0]) begin
          coeffs_133 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_134 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h86 == rs2[9:0]) begin
          coeffs_134 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_135 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h87 == rs2[9:0]) begin
          coeffs_135 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_136 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h88 == rs2[9:0]) begin
          coeffs_136 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_137 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h89 == rs2[9:0]) begin
          coeffs_137 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_138 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h8a == rs2[9:0]) begin
          coeffs_138 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_139 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h8b == rs2[9:0]) begin
          coeffs_139 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_140 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h8c == rs2[9:0]) begin
          coeffs_140 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_141 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h8d == rs2[9:0]) begin
          coeffs_141 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_142 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h8e == rs2[9:0]) begin
          coeffs_142 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_143 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h8f == rs2[9:0]) begin
          coeffs_143 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_144 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h90 == rs2[9:0]) begin
          coeffs_144 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_145 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h91 == rs2[9:0]) begin
          coeffs_145 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_146 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h92 == rs2[9:0]) begin
          coeffs_146 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_147 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h93 == rs2[9:0]) begin
          coeffs_147 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_148 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h94 == rs2[9:0]) begin
          coeffs_148 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_149 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h95 == rs2[9:0]) begin
          coeffs_149 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_150 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h96 == rs2[9:0]) begin
          coeffs_150 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_151 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h97 == rs2[9:0]) begin
          coeffs_151 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_152 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h98 == rs2[9:0]) begin
          coeffs_152 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_153 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h99 == rs2[9:0]) begin
          coeffs_153 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_154 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h9a == rs2[9:0]) begin
          coeffs_154 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_155 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h9b == rs2[9:0]) begin
          coeffs_155 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_156 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h9c == rs2[9:0]) begin
          coeffs_156 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_157 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h9d == rs2[9:0]) begin
          coeffs_157 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_158 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h9e == rs2[9:0]) begin
          coeffs_158 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_159 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h9f == rs2[9:0]) begin
          coeffs_159 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_160 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha0 == rs2[9:0]) begin
          coeffs_160 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_161 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha1 == rs2[9:0]) begin
          coeffs_161 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_162 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha2 == rs2[9:0]) begin
          coeffs_162 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_163 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha3 == rs2[9:0]) begin
          coeffs_163 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_164 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha4 == rs2[9:0]) begin
          coeffs_164 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_165 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha5 == rs2[9:0]) begin
          coeffs_165 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_166 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha6 == rs2[9:0]) begin
          coeffs_166 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_167 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha7 == rs2[9:0]) begin
          coeffs_167 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_168 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha8 == rs2[9:0]) begin
          coeffs_168 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_169 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'ha9 == rs2[9:0]) begin
          coeffs_169 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_170 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'haa == rs2[9:0]) begin
          coeffs_170 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_171 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hab == rs2[9:0]) begin
          coeffs_171 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_172 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hac == rs2[9:0]) begin
          coeffs_172 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_173 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'had == rs2[9:0]) begin
          coeffs_173 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_174 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hae == rs2[9:0]) begin
          coeffs_174 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_175 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'haf == rs2[9:0]) begin
          coeffs_175 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_176 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb0 == rs2[9:0]) begin
          coeffs_176 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_177 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb1 == rs2[9:0]) begin
          coeffs_177 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_178 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb2 == rs2[9:0]) begin
          coeffs_178 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_179 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb3 == rs2[9:0]) begin
          coeffs_179 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_180 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb4 == rs2[9:0]) begin
          coeffs_180 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_181 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb5 == rs2[9:0]) begin
          coeffs_181 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_182 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb6 == rs2[9:0]) begin
          coeffs_182 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_183 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb7 == rs2[9:0]) begin
          coeffs_183 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_184 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb8 == rs2[9:0]) begin
          coeffs_184 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_185 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hb9 == rs2[9:0]) begin
          coeffs_185 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_186 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hba == rs2[9:0]) begin
          coeffs_186 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_187 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hbb == rs2[9:0]) begin
          coeffs_187 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_188 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hbc == rs2[9:0]) begin
          coeffs_188 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_189 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hbd == rs2[9:0]) begin
          coeffs_189 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_190 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hbe == rs2[9:0]) begin
          coeffs_190 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_191 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hbf == rs2[9:0]) begin
          coeffs_191 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_192 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc0 == rs2[9:0]) begin
          coeffs_192 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_193 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc1 == rs2[9:0]) begin
          coeffs_193 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_194 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc2 == rs2[9:0]) begin
          coeffs_194 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_195 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc3 == rs2[9:0]) begin
          coeffs_195 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_196 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc4 == rs2[9:0]) begin
          coeffs_196 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_197 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc5 == rs2[9:0]) begin
          coeffs_197 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_198 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc6 == rs2[9:0]) begin
          coeffs_198 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_199 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc7 == rs2[9:0]) begin
          coeffs_199 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_200 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc8 == rs2[9:0]) begin
          coeffs_200 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_201 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hc9 == rs2[9:0]) begin
          coeffs_201 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_202 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hca == rs2[9:0]) begin
          coeffs_202 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_203 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hcb == rs2[9:0]) begin
          coeffs_203 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_204 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hcc == rs2[9:0]) begin
          coeffs_204 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_205 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hcd == rs2[9:0]) begin
          coeffs_205 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_206 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hce == rs2[9:0]) begin
          coeffs_206 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_207 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hcf == rs2[9:0]) begin
          coeffs_207 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_208 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd0 == rs2[9:0]) begin
          coeffs_208 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_209 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd1 == rs2[9:0]) begin
          coeffs_209 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_210 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd2 == rs2[9:0]) begin
          coeffs_210 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_211 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd3 == rs2[9:0]) begin
          coeffs_211 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_212 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd4 == rs2[9:0]) begin
          coeffs_212 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_213 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd5 == rs2[9:0]) begin
          coeffs_213 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_214 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd6 == rs2[9:0]) begin
          coeffs_214 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_215 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd7 == rs2[9:0]) begin
          coeffs_215 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_216 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd8 == rs2[9:0]) begin
          coeffs_216 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_217 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hd9 == rs2[9:0]) begin
          coeffs_217 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_218 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hda == rs2[9:0]) begin
          coeffs_218 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_219 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hdb == rs2[9:0]) begin
          coeffs_219 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_220 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hdc == rs2[9:0]) begin
          coeffs_220 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_221 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hdd == rs2[9:0]) begin
          coeffs_221 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_222 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hde == rs2[9:0]) begin
          coeffs_222 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_223 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hdf == rs2[9:0]) begin
          coeffs_223 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_224 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he0 == rs2[9:0]) begin
          coeffs_224 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_225 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he1 == rs2[9:0]) begin
          coeffs_225 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_226 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he2 == rs2[9:0]) begin
          coeffs_226 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_227 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he3 == rs2[9:0]) begin
          coeffs_227 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_228 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he4 == rs2[9:0]) begin
          coeffs_228 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_229 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he5 == rs2[9:0]) begin
          coeffs_229 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_230 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he6 == rs2[9:0]) begin
          coeffs_230 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_231 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he7 == rs2[9:0]) begin
          coeffs_231 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_232 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he8 == rs2[9:0]) begin
          coeffs_232 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_233 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'he9 == rs2[9:0]) begin
          coeffs_233 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_234 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hea == rs2[9:0]) begin
          coeffs_234 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_235 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'heb == rs2[9:0]) begin
          coeffs_235 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_236 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hec == rs2[9:0]) begin
          coeffs_236 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_237 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hed == rs2[9:0]) begin
          coeffs_237 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_238 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hee == rs2[9:0]) begin
          coeffs_238 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_239 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hef == rs2[9:0]) begin
          coeffs_239 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_240 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf0 == rs2[9:0]) begin
          coeffs_240 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_241 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf1 == rs2[9:0]) begin
          coeffs_241 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_242 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf2 == rs2[9:0]) begin
          coeffs_242 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_243 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf3 == rs2[9:0]) begin
          coeffs_243 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_244 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf4 == rs2[9:0]) begin
          coeffs_244 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_245 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf5 == rs2[9:0]) begin
          coeffs_245 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_246 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf6 == rs2[9:0]) begin
          coeffs_246 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_247 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf7 == rs2[9:0]) begin
          coeffs_247 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_248 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf8 == rs2[9:0]) begin
          coeffs_248 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_249 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hf9 == rs2[9:0]) begin
          coeffs_249 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_250 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hfa == rs2[9:0]) begin
          coeffs_250 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_251 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hfb == rs2[9:0]) begin
          coeffs_251 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_252 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hfc == rs2[9:0]) begin
          coeffs_252 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_253 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hfd == rs2[9:0]) begin
          coeffs_253 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_254 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hfe == rs2[9:0]) begin
          coeffs_254 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_255 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'hff == rs2[9:0]) begin
          coeffs_255 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_256 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h100 == rs2[9:0]) begin
          coeffs_256 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_257 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h101 == rs2[9:0]) begin
          coeffs_257 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_258 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h102 == rs2[9:0]) begin
          coeffs_258 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_259 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h103 == rs2[9:0]) begin
          coeffs_259 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_260 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h104 == rs2[9:0]) begin
          coeffs_260 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_261 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h105 == rs2[9:0]) begin
          coeffs_261 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_262 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h106 == rs2[9:0]) begin
          coeffs_262 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_263 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h107 == rs2[9:0]) begin
          coeffs_263 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_264 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h108 == rs2[9:0]) begin
          coeffs_264 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_265 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h109 == rs2[9:0]) begin
          coeffs_265 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_266 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h10a == rs2[9:0]) begin
          coeffs_266 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_267 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h10b == rs2[9:0]) begin
          coeffs_267 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_268 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h10c == rs2[9:0]) begin
          coeffs_268 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_269 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h10d == rs2[9:0]) begin
          coeffs_269 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_270 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h10e == rs2[9:0]) begin
          coeffs_270 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_271 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h10f == rs2[9:0]) begin
          coeffs_271 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_272 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h110 == rs2[9:0]) begin
          coeffs_272 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_273 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h111 == rs2[9:0]) begin
          coeffs_273 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_274 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h112 == rs2[9:0]) begin
          coeffs_274 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_275 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h113 == rs2[9:0]) begin
          coeffs_275 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_276 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h114 == rs2[9:0]) begin
          coeffs_276 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_277 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h115 == rs2[9:0]) begin
          coeffs_277 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_278 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h116 == rs2[9:0]) begin
          coeffs_278 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_279 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h117 == rs2[9:0]) begin
          coeffs_279 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_280 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h118 == rs2[9:0]) begin
          coeffs_280 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_281 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h119 == rs2[9:0]) begin
          coeffs_281 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_282 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h11a == rs2[9:0]) begin
          coeffs_282 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_283 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h11b == rs2[9:0]) begin
          coeffs_283 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_284 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h11c == rs2[9:0]) begin
          coeffs_284 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_285 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h11d == rs2[9:0]) begin
          coeffs_285 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_286 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h11e == rs2[9:0]) begin
          coeffs_286 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_287 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h11f == rs2[9:0]) begin
          coeffs_287 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_288 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h120 == rs2[9:0]) begin
          coeffs_288 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_289 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h121 == rs2[9:0]) begin
          coeffs_289 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_290 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h122 == rs2[9:0]) begin
          coeffs_290 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_291 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h123 == rs2[9:0]) begin
          coeffs_291 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_292 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h124 == rs2[9:0]) begin
          coeffs_292 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_293 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h125 == rs2[9:0]) begin
          coeffs_293 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_294 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h126 == rs2[9:0]) begin
          coeffs_294 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_295 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h127 == rs2[9:0]) begin
          coeffs_295 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_296 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h128 == rs2[9:0]) begin
          coeffs_296 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_297 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h129 == rs2[9:0]) begin
          coeffs_297 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_298 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h12a == rs2[9:0]) begin
          coeffs_298 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_299 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h12b == rs2[9:0]) begin
          coeffs_299 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_300 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h12c == rs2[9:0]) begin
          coeffs_300 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_301 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h12d == rs2[9:0]) begin
          coeffs_301 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_302 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h12e == rs2[9:0]) begin
          coeffs_302 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_303 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h12f == rs2[9:0]) begin
          coeffs_303 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_304 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h130 == rs2[9:0]) begin
          coeffs_304 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_305 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h131 == rs2[9:0]) begin
          coeffs_305 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_306 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h132 == rs2[9:0]) begin
          coeffs_306 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_307 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h133 == rs2[9:0]) begin
          coeffs_307 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_308 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h134 == rs2[9:0]) begin
          coeffs_308 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_309 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h135 == rs2[9:0]) begin
          coeffs_309 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_310 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h136 == rs2[9:0]) begin
          coeffs_310 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_311 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h137 == rs2[9:0]) begin
          coeffs_311 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_312 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h138 == rs2[9:0]) begin
          coeffs_312 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_313 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h139 == rs2[9:0]) begin
          coeffs_313 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_314 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h13a == rs2[9:0]) begin
          coeffs_314 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_315 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h13b == rs2[9:0]) begin
          coeffs_315 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_316 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h13c == rs2[9:0]) begin
          coeffs_316 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_317 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h13d == rs2[9:0]) begin
          coeffs_317 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_318 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h13e == rs2[9:0]) begin
          coeffs_318 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_319 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h13f == rs2[9:0]) begin
          coeffs_319 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_320 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h140 == rs2[9:0]) begin
          coeffs_320 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_321 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h141 == rs2[9:0]) begin
          coeffs_321 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_322 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h142 == rs2[9:0]) begin
          coeffs_322 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_323 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h143 == rs2[9:0]) begin
          coeffs_323 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_324 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h144 == rs2[9:0]) begin
          coeffs_324 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_325 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h145 == rs2[9:0]) begin
          coeffs_325 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_326 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h146 == rs2[9:0]) begin
          coeffs_326 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_327 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h147 == rs2[9:0]) begin
          coeffs_327 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_328 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h148 == rs2[9:0]) begin
          coeffs_328 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_329 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h149 == rs2[9:0]) begin
          coeffs_329 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_330 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h14a == rs2[9:0]) begin
          coeffs_330 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_331 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h14b == rs2[9:0]) begin
          coeffs_331 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_332 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h14c == rs2[9:0]) begin
          coeffs_332 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_333 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h14d == rs2[9:0]) begin
          coeffs_333 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_334 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h14e == rs2[9:0]) begin
          coeffs_334 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_335 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h14f == rs2[9:0]) begin
          coeffs_335 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_336 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h150 == rs2[9:0]) begin
          coeffs_336 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_337 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h151 == rs2[9:0]) begin
          coeffs_337 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_338 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h152 == rs2[9:0]) begin
          coeffs_338 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_339 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h153 == rs2[9:0]) begin
          coeffs_339 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_340 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h154 == rs2[9:0]) begin
          coeffs_340 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_341 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h155 == rs2[9:0]) begin
          coeffs_341 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_342 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h156 == rs2[9:0]) begin
          coeffs_342 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_343 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h157 == rs2[9:0]) begin
          coeffs_343 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_344 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h158 == rs2[9:0]) begin
          coeffs_344 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_345 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h159 == rs2[9:0]) begin
          coeffs_345 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_346 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h15a == rs2[9:0]) begin
          coeffs_346 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_347 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h15b == rs2[9:0]) begin
          coeffs_347 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_348 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h15c == rs2[9:0]) begin
          coeffs_348 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_349 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h15d == rs2[9:0]) begin
          coeffs_349 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_350 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h15e == rs2[9:0]) begin
          coeffs_350 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_351 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h15f == rs2[9:0]) begin
          coeffs_351 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_352 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h160 == rs2[9:0]) begin
          coeffs_352 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_353 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h161 == rs2[9:0]) begin
          coeffs_353 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_354 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h162 == rs2[9:0]) begin
          coeffs_354 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_355 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h163 == rs2[9:0]) begin
          coeffs_355 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_356 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h164 == rs2[9:0]) begin
          coeffs_356 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_357 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h165 == rs2[9:0]) begin
          coeffs_357 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_358 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h166 == rs2[9:0]) begin
          coeffs_358 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_359 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h167 == rs2[9:0]) begin
          coeffs_359 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_360 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h168 == rs2[9:0]) begin
          coeffs_360 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_361 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h169 == rs2[9:0]) begin
          coeffs_361 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_362 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h16a == rs2[9:0]) begin
          coeffs_362 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_363 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h16b == rs2[9:0]) begin
          coeffs_363 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_364 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h16c == rs2[9:0]) begin
          coeffs_364 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_365 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h16d == rs2[9:0]) begin
          coeffs_365 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_366 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h16e == rs2[9:0]) begin
          coeffs_366 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_367 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h16f == rs2[9:0]) begin
          coeffs_367 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_368 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h170 == rs2[9:0]) begin
          coeffs_368 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_369 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h171 == rs2[9:0]) begin
          coeffs_369 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_370 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h172 == rs2[9:0]) begin
          coeffs_370 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_371 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h173 == rs2[9:0]) begin
          coeffs_371 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_372 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h174 == rs2[9:0]) begin
          coeffs_372 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_373 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h175 == rs2[9:0]) begin
          coeffs_373 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_374 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h176 == rs2[9:0]) begin
          coeffs_374 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_375 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h177 == rs2[9:0]) begin
          coeffs_375 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_376 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h178 == rs2[9:0]) begin
          coeffs_376 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_377 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h179 == rs2[9:0]) begin
          coeffs_377 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_378 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h17a == rs2[9:0]) begin
          coeffs_378 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_379 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h17b == rs2[9:0]) begin
          coeffs_379 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_380 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h17c == rs2[9:0]) begin
          coeffs_380 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_381 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h17d == rs2[9:0]) begin
          coeffs_381 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_382 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h17e == rs2[9:0]) begin
          coeffs_382 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_383 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h17f == rs2[9:0]) begin
          coeffs_383 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_384 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h180 == rs2[9:0]) begin
          coeffs_384 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_385 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h181 == rs2[9:0]) begin
          coeffs_385 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_386 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h182 == rs2[9:0]) begin
          coeffs_386 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_387 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h183 == rs2[9:0]) begin
          coeffs_387 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_388 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h184 == rs2[9:0]) begin
          coeffs_388 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_389 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h185 == rs2[9:0]) begin
          coeffs_389 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_390 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h186 == rs2[9:0]) begin
          coeffs_390 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_391 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h187 == rs2[9:0]) begin
          coeffs_391 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_392 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h188 == rs2[9:0]) begin
          coeffs_392 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_393 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h189 == rs2[9:0]) begin
          coeffs_393 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_394 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h18a == rs2[9:0]) begin
          coeffs_394 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_395 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h18b == rs2[9:0]) begin
          coeffs_395 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_396 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h18c == rs2[9:0]) begin
          coeffs_396 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_397 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h18d == rs2[9:0]) begin
          coeffs_397 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_398 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h18e == rs2[9:0]) begin
          coeffs_398 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_399 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h18f == rs2[9:0]) begin
          coeffs_399 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_400 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h190 == rs2[9:0]) begin
          coeffs_400 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_401 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h191 == rs2[9:0]) begin
          coeffs_401 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_402 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h192 == rs2[9:0]) begin
          coeffs_402 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_403 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h193 == rs2[9:0]) begin
          coeffs_403 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_404 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h194 == rs2[9:0]) begin
          coeffs_404 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_405 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h195 == rs2[9:0]) begin
          coeffs_405 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_406 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h196 == rs2[9:0]) begin
          coeffs_406 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_407 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h197 == rs2[9:0]) begin
          coeffs_407 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_408 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h198 == rs2[9:0]) begin
          coeffs_408 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_409 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h199 == rs2[9:0]) begin
          coeffs_409 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_410 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h19a == rs2[9:0]) begin
          coeffs_410 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_411 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h19b == rs2[9:0]) begin
          coeffs_411 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_412 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h19c == rs2[9:0]) begin
          coeffs_412 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_413 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h19d == rs2[9:0]) begin
          coeffs_413 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_414 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h19e == rs2[9:0]) begin
          coeffs_414 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_415 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h19f == rs2[9:0]) begin
          coeffs_415 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_416 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a0 == rs2[9:0]) begin
          coeffs_416 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_417 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a1 == rs2[9:0]) begin
          coeffs_417 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_418 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a2 == rs2[9:0]) begin
          coeffs_418 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_419 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a3 == rs2[9:0]) begin
          coeffs_419 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_420 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a4 == rs2[9:0]) begin
          coeffs_420 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_421 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a5 == rs2[9:0]) begin
          coeffs_421 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_422 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a6 == rs2[9:0]) begin
          coeffs_422 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_423 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a7 == rs2[9:0]) begin
          coeffs_423 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_424 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a8 == rs2[9:0]) begin
          coeffs_424 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_425 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1a9 == rs2[9:0]) begin
          coeffs_425 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_426 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1aa == rs2[9:0]) begin
          coeffs_426 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_427 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ab == rs2[9:0]) begin
          coeffs_427 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_428 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ac == rs2[9:0]) begin
          coeffs_428 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_429 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ad == rs2[9:0]) begin
          coeffs_429 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_430 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ae == rs2[9:0]) begin
          coeffs_430 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_431 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1af == rs2[9:0]) begin
          coeffs_431 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_432 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b0 == rs2[9:0]) begin
          coeffs_432 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_433 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b1 == rs2[9:0]) begin
          coeffs_433 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_434 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b2 == rs2[9:0]) begin
          coeffs_434 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_435 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b3 == rs2[9:0]) begin
          coeffs_435 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_436 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b4 == rs2[9:0]) begin
          coeffs_436 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_437 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b5 == rs2[9:0]) begin
          coeffs_437 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_438 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b6 == rs2[9:0]) begin
          coeffs_438 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_439 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b7 == rs2[9:0]) begin
          coeffs_439 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_440 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b8 == rs2[9:0]) begin
          coeffs_440 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_441 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1b9 == rs2[9:0]) begin
          coeffs_441 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_442 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ba == rs2[9:0]) begin
          coeffs_442 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_443 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1bb == rs2[9:0]) begin
          coeffs_443 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_444 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1bc == rs2[9:0]) begin
          coeffs_444 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_445 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1bd == rs2[9:0]) begin
          coeffs_445 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_446 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1be == rs2[9:0]) begin
          coeffs_446 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_447 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1bf == rs2[9:0]) begin
          coeffs_447 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_448 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c0 == rs2[9:0]) begin
          coeffs_448 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_449 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c1 == rs2[9:0]) begin
          coeffs_449 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_450 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c2 == rs2[9:0]) begin
          coeffs_450 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_451 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c3 == rs2[9:0]) begin
          coeffs_451 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_452 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c4 == rs2[9:0]) begin
          coeffs_452 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_453 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c5 == rs2[9:0]) begin
          coeffs_453 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_454 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c6 == rs2[9:0]) begin
          coeffs_454 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_455 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c7 == rs2[9:0]) begin
          coeffs_455 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_456 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c8 == rs2[9:0]) begin
          coeffs_456 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_457 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1c9 == rs2[9:0]) begin
          coeffs_457 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_458 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ca == rs2[9:0]) begin
          coeffs_458 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_459 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1cb == rs2[9:0]) begin
          coeffs_459 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_460 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1cc == rs2[9:0]) begin
          coeffs_460 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_461 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1cd == rs2[9:0]) begin
          coeffs_461 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_462 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ce == rs2[9:0]) begin
          coeffs_462 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_463 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1cf == rs2[9:0]) begin
          coeffs_463 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_464 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d0 == rs2[9:0]) begin
          coeffs_464 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_465 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d1 == rs2[9:0]) begin
          coeffs_465 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_466 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d2 == rs2[9:0]) begin
          coeffs_466 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_467 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d3 == rs2[9:0]) begin
          coeffs_467 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_468 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d4 == rs2[9:0]) begin
          coeffs_468 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_469 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d5 == rs2[9:0]) begin
          coeffs_469 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_470 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d6 == rs2[9:0]) begin
          coeffs_470 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_471 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d7 == rs2[9:0]) begin
          coeffs_471 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_472 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d8 == rs2[9:0]) begin
          coeffs_472 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_473 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1d9 == rs2[9:0]) begin
          coeffs_473 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_474 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1da == rs2[9:0]) begin
          coeffs_474 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_475 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1db == rs2[9:0]) begin
          coeffs_475 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_476 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1dc == rs2[9:0]) begin
          coeffs_476 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_477 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1dd == rs2[9:0]) begin
          coeffs_477 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_478 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1de == rs2[9:0]) begin
          coeffs_478 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_479 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1df == rs2[9:0]) begin
          coeffs_479 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_480 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e0 == rs2[9:0]) begin
          coeffs_480 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_481 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e1 == rs2[9:0]) begin
          coeffs_481 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_482 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e2 == rs2[9:0]) begin
          coeffs_482 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_483 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e3 == rs2[9:0]) begin
          coeffs_483 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_484 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e4 == rs2[9:0]) begin
          coeffs_484 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_485 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e5 == rs2[9:0]) begin
          coeffs_485 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_486 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e6 == rs2[9:0]) begin
          coeffs_486 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_487 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e7 == rs2[9:0]) begin
          coeffs_487 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_488 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e8 == rs2[9:0]) begin
          coeffs_488 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_489 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1e9 == rs2[9:0]) begin
          coeffs_489 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_490 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ea == rs2[9:0]) begin
          coeffs_490 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_491 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1eb == rs2[9:0]) begin
          coeffs_491 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_492 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ec == rs2[9:0]) begin
          coeffs_492 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_493 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ed == rs2[9:0]) begin
          coeffs_493 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_494 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ee == rs2[9:0]) begin
          coeffs_494 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_495 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ef == rs2[9:0]) begin
          coeffs_495 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_496 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f0 == rs2[9:0]) begin
          coeffs_496 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_497 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f1 == rs2[9:0]) begin
          coeffs_497 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_498 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f2 == rs2[9:0]) begin
          coeffs_498 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_499 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f3 == rs2[9:0]) begin
          coeffs_499 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_500 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f4 == rs2[9:0]) begin
          coeffs_500 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_501 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f5 == rs2[9:0]) begin
          coeffs_501 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_502 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f6 == rs2[9:0]) begin
          coeffs_502 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_503 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f7 == rs2[9:0]) begin
          coeffs_503 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_504 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f8 == rs2[9:0]) begin
          coeffs_504 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_505 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1f9 == rs2[9:0]) begin
          coeffs_505 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_506 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1fa == rs2[9:0]) begin
          coeffs_506 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_507 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1fb == rs2[9:0]) begin
          coeffs_507 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_508 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1fc == rs2[9:0]) begin
          coeffs_508 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_509 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1fd == rs2[9:0]) begin
          coeffs_509 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_510 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1fe == rs2[9:0]) begin
          coeffs_510 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_511 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h1ff == rs2[9:0]) begin
          coeffs_511 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_512 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h200 == rs2[9:0]) begin
          coeffs_512 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_513 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h201 == rs2[9:0]) begin
          coeffs_513 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_514 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h202 == rs2[9:0]) begin
          coeffs_514 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_515 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h203 == rs2[9:0]) begin
          coeffs_515 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_516 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h204 == rs2[9:0]) begin
          coeffs_516 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_517 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h205 == rs2[9:0]) begin
          coeffs_517 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_518 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h206 == rs2[9:0]) begin
          coeffs_518 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_519 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h207 == rs2[9:0]) begin
          coeffs_519 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_520 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h208 == rs2[9:0]) begin
          coeffs_520 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_521 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h209 == rs2[9:0]) begin
          coeffs_521 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_522 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h20a == rs2[9:0]) begin
          coeffs_522 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_523 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h20b == rs2[9:0]) begin
          coeffs_523 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_524 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h20c == rs2[9:0]) begin
          coeffs_524 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_525 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h20d == rs2[9:0]) begin
          coeffs_525 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_526 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h20e == rs2[9:0]) begin
          coeffs_526 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_527 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h20f == rs2[9:0]) begin
          coeffs_527 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_528 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h210 == rs2[9:0]) begin
          coeffs_528 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_529 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h211 == rs2[9:0]) begin
          coeffs_529 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_530 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h212 == rs2[9:0]) begin
          coeffs_530 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_531 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h213 == rs2[9:0]) begin
          coeffs_531 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_532 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h214 == rs2[9:0]) begin
          coeffs_532 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_533 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h215 == rs2[9:0]) begin
          coeffs_533 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_534 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h216 == rs2[9:0]) begin
          coeffs_534 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_535 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h217 == rs2[9:0]) begin
          coeffs_535 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_536 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h218 == rs2[9:0]) begin
          coeffs_536 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_537 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h219 == rs2[9:0]) begin
          coeffs_537 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_538 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h21a == rs2[9:0]) begin
          coeffs_538 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_539 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h21b == rs2[9:0]) begin
          coeffs_539 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_540 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h21c == rs2[9:0]) begin
          coeffs_540 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_541 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h21d == rs2[9:0]) begin
          coeffs_541 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_542 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h21e == rs2[9:0]) begin
          coeffs_542 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_543 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h21f == rs2[9:0]) begin
          coeffs_543 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_544 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h220 == rs2[9:0]) begin
          coeffs_544 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_545 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h221 == rs2[9:0]) begin
          coeffs_545 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_546 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h222 == rs2[9:0]) begin
          coeffs_546 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_547 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h223 == rs2[9:0]) begin
          coeffs_547 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_548 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h224 == rs2[9:0]) begin
          coeffs_548 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_549 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h225 == rs2[9:0]) begin
          coeffs_549 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_550 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h226 == rs2[9:0]) begin
          coeffs_550 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_551 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h227 == rs2[9:0]) begin
          coeffs_551 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_552 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h228 == rs2[9:0]) begin
          coeffs_552 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_553 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h229 == rs2[9:0]) begin
          coeffs_553 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_554 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h22a == rs2[9:0]) begin
          coeffs_554 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_555 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h22b == rs2[9:0]) begin
          coeffs_555 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_556 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h22c == rs2[9:0]) begin
          coeffs_556 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_557 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h22d == rs2[9:0]) begin
          coeffs_557 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_558 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h22e == rs2[9:0]) begin
          coeffs_558 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_559 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h22f == rs2[9:0]) begin
          coeffs_559 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_560 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h230 == rs2[9:0]) begin
          coeffs_560 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_561 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h231 == rs2[9:0]) begin
          coeffs_561 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_562 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h232 == rs2[9:0]) begin
          coeffs_562 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_563 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h233 == rs2[9:0]) begin
          coeffs_563 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_564 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h234 == rs2[9:0]) begin
          coeffs_564 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_565 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h235 == rs2[9:0]) begin
          coeffs_565 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_566 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h236 == rs2[9:0]) begin
          coeffs_566 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_567 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h237 == rs2[9:0]) begin
          coeffs_567 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_568 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h238 == rs2[9:0]) begin
          coeffs_568 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_569 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h239 == rs2[9:0]) begin
          coeffs_569 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_570 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h23a == rs2[9:0]) begin
          coeffs_570 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_571 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h23b == rs2[9:0]) begin
          coeffs_571 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_572 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h23c == rs2[9:0]) begin
          coeffs_572 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_573 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h23d == rs2[9:0]) begin
          coeffs_573 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_574 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h23e == rs2[9:0]) begin
          coeffs_574 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_575 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h23f == rs2[9:0]) begin
          coeffs_575 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_576 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h240 == rs2[9:0]) begin
          coeffs_576 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_577 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h241 == rs2[9:0]) begin
          coeffs_577 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_578 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h242 == rs2[9:0]) begin
          coeffs_578 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_579 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h243 == rs2[9:0]) begin
          coeffs_579 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_580 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h244 == rs2[9:0]) begin
          coeffs_580 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_581 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h245 == rs2[9:0]) begin
          coeffs_581 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_582 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h246 == rs2[9:0]) begin
          coeffs_582 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_583 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h247 == rs2[9:0]) begin
          coeffs_583 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_584 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h248 == rs2[9:0]) begin
          coeffs_584 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_585 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h249 == rs2[9:0]) begin
          coeffs_585 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_586 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h24a == rs2[9:0]) begin
          coeffs_586 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_587 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h24b == rs2[9:0]) begin
          coeffs_587 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_588 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h24c == rs2[9:0]) begin
          coeffs_588 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_589 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h24d == rs2[9:0]) begin
          coeffs_589 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_590 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h24e == rs2[9:0]) begin
          coeffs_590 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_591 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h24f == rs2[9:0]) begin
          coeffs_591 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_592 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h250 == rs2[9:0]) begin
          coeffs_592 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_593 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h251 == rs2[9:0]) begin
          coeffs_593 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_594 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h252 == rs2[9:0]) begin
          coeffs_594 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_595 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h253 == rs2[9:0]) begin
          coeffs_595 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_596 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h254 == rs2[9:0]) begin
          coeffs_596 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_597 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h255 == rs2[9:0]) begin
          coeffs_597 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_598 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h256 == rs2[9:0]) begin
          coeffs_598 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_599 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h257 == rs2[9:0]) begin
          coeffs_599 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_600 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h258 == rs2[9:0]) begin
          coeffs_600 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_601 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h259 == rs2[9:0]) begin
          coeffs_601 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_602 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h25a == rs2[9:0]) begin
          coeffs_602 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_603 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h25b == rs2[9:0]) begin
          coeffs_603 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_604 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h25c == rs2[9:0]) begin
          coeffs_604 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_605 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h25d == rs2[9:0]) begin
          coeffs_605 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_606 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h25e == rs2[9:0]) begin
          coeffs_606 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_607 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h25f == rs2[9:0]) begin
          coeffs_607 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_608 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h260 == rs2[9:0]) begin
          coeffs_608 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_609 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h261 == rs2[9:0]) begin
          coeffs_609 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_610 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h262 == rs2[9:0]) begin
          coeffs_610 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_611 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h263 == rs2[9:0]) begin
          coeffs_611 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_612 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h264 == rs2[9:0]) begin
          coeffs_612 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_613 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h265 == rs2[9:0]) begin
          coeffs_613 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_614 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h266 == rs2[9:0]) begin
          coeffs_614 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_615 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h267 == rs2[9:0]) begin
          coeffs_615 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_616 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h268 == rs2[9:0]) begin
          coeffs_616 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_617 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h269 == rs2[9:0]) begin
          coeffs_617 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_618 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h26a == rs2[9:0]) begin
          coeffs_618 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_619 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h26b == rs2[9:0]) begin
          coeffs_619 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_620 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h26c == rs2[9:0]) begin
          coeffs_620 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_621 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h26d == rs2[9:0]) begin
          coeffs_621 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_622 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h26e == rs2[9:0]) begin
          coeffs_622 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_623 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h26f == rs2[9:0]) begin
          coeffs_623 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_624 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h270 == rs2[9:0]) begin
          coeffs_624 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_625 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h271 == rs2[9:0]) begin
          coeffs_625 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_626 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h272 == rs2[9:0]) begin
          coeffs_626 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_627 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h273 == rs2[9:0]) begin
          coeffs_627 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_628 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h274 == rs2[9:0]) begin
          coeffs_628 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_629 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h275 == rs2[9:0]) begin
          coeffs_629 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_630 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h276 == rs2[9:0]) begin
          coeffs_630 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_631 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h277 == rs2[9:0]) begin
          coeffs_631 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_632 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h278 == rs2[9:0]) begin
          coeffs_632 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_633 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h279 == rs2[9:0]) begin
          coeffs_633 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_634 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h27a == rs2[9:0]) begin
          coeffs_634 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_635 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h27b == rs2[9:0]) begin
          coeffs_635 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_636 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h27c == rs2[9:0]) begin
          coeffs_636 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_637 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h27d == rs2[9:0]) begin
          coeffs_637 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_638 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h27e == rs2[9:0]) begin
          coeffs_638 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_639 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h27f == rs2[9:0]) begin
          coeffs_639 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_640 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h280 == rs2[9:0]) begin
          coeffs_640 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_641 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h281 == rs2[9:0]) begin
          coeffs_641 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_642 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h282 == rs2[9:0]) begin
          coeffs_642 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_643 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h283 == rs2[9:0]) begin
          coeffs_643 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_644 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h284 == rs2[9:0]) begin
          coeffs_644 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_645 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h285 == rs2[9:0]) begin
          coeffs_645 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_646 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h286 == rs2[9:0]) begin
          coeffs_646 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_647 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h287 == rs2[9:0]) begin
          coeffs_647 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_648 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h288 == rs2[9:0]) begin
          coeffs_648 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_649 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h289 == rs2[9:0]) begin
          coeffs_649 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_650 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h28a == rs2[9:0]) begin
          coeffs_650 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_651 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h28b == rs2[9:0]) begin
          coeffs_651 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_652 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h28c == rs2[9:0]) begin
          coeffs_652 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_653 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h28d == rs2[9:0]) begin
          coeffs_653 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_654 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h28e == rs2[9:0]) begin
          coeffs_654 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_655 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h28f == rs2[9:0]) begin
          coeffs_655 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_656 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h290 == rs2[9:0]) begin
          coeffs_656 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_657 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h291 == rs2[9:0]) begin
          coeffs_657 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_658 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h292 == rs2[9:0]) begin
          coeffs_658 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_659 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h293 == rs2[9:0]) begin
          coeffs_659 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_660 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h294 == rs2[9:0]) begin
          coeffs_660 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_661 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h295 == rs2[9:0]) begin
          coeffs_661 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_662 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h296 == rs2[9:0]) begin
          coeffs_662 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_663 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h297 == rs2[9:0]) begin
          coeffs_663 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_664 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h298 == rs2[9:0]) begin
          coeffs_664 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_665 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h299 == rs2[9:0]) begin
          coeffs_665 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_666 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h29a == rs2[9:0]) begin
          coeffs_666 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_667 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h29b == rs2[9:0]) begin
          coeffs_667 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_668 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h29c == rs2[9:0]) begin
          coeffs_668 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_669 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h29d == rs2[9:0]) begin
          coeffs_669 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_670 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h29e == rs2[9:0]) begin
          coeffs_670 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_671 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h29f == rs2[9:0]) begin
          coeffs_671 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_672 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a0 == rs2[9:0]) begin
          coeffs_672 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_673 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a1 == rs2[9:0]) begin
          coeffs_673 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_674 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a2 == rs2[9:0]) begin
          coeffs_674 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_675 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a3 == rs2[9:0]) begin
          coeffs_675 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_676 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a4 == rs2[9:0]) begin
          coeffs_676 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_677 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a5 == rs2[9:0]) begin
          coeffs_677 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_678 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a6 == rs2[9:0]) begin
          coeffs_678 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_679 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a7 == rs2[9:0]) begin
          coeffs_679 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_680 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a8 == rs2[9:0]) begin
          coeffs_680 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_681 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2a9 == rs2[9:0]) begin
          coeffs_681 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_682 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2aa == rs2[9:0]) begin
          coeffs_682 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_683 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ab == rs2[9:0]) begin
          coeffs_683 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_684 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ac == rs2[9:0]) begin
          coeffs_684 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_685 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ad == rs2[9:0]) begin
          coeffs_685 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_686 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ae == rs2[9:0]) begin
          coeffs_686 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_687 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2af == rs2[9:0]) begin
          coeffs_687 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_688 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b0 == rs2[9:0]) begin
          coeffs_688 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_689 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b1 == rs2[9:0]) begin
          coeffs_689 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_690 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b2 == rs2[9:0]) begin
          coeffs_690 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_691 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b3 == rs2[9:0]) begin
          coeffs_691 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_692 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b4 == rs2[9:0]) begin
          coeffs_692 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_693 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b5 == rs2[9:0]) begin
          coeffs_693 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_694 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b6 == rs2[9:0]) begin
          coeffs_694 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_695 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b7 == rs2[9:0]) begin
          coeffs_695 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_696 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b8 == rs2[9:0]) begin
          coeffs_696 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_697 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2b9 == rs2[9:0]) begin
          coeffs_697 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_698 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ba == rs2[9:0]) begin
          coeffs_698 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_699 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2bb == rs2[9:0]) begin
          coeffs_699 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_700 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2bc == rs2[9:0]) begin
          coeffs_700 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_701 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2bd == rs2[9:0]) begin
          coeffs_701 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_702 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2be == rs2[9:0]) begin
          coeffs_702 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_703 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2bf == rs2[9:0]) begin
          coeffs_703 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_704 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c0 == rs2[9:0]) begin
          coeffs_704 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_705 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c1 == rs2[9:0]) begin
          coeffs_705 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_706 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c2 == rs2[9:0]) begin
          coeffs_706 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_707 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c3 == rs2[9:0]) begin
          coeffs_707 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_708 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c4 == rs2[9:0]) begin
          coeffs_708 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_709 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c5 == rs2[9:0]) begin
          coeffs_709 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_710 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c6 == rs2[9:0]) begin
          coeffs_710 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_711 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c7 == rs2[9:0]) begin
          coeffs_711 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_712 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c8 == rs2[9:0]) begin
          coeffs_712 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_713 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2c9 == rs2[9:0]) begin
          coeffs_713 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_714 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ca == rs2[9:0]) begin
          coeffs_714 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_715 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2cb == rs2[9:0]) begin
          coeffs_715 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_716 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2cc == rs2[9:0]) begin
          coeffs_716 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_717 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2cd == rs2[9:0]) begin
          coeffs_717 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_718 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ce == rs2[9:0]) begin
          coeffs_718 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_719 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2cf == rs2[9:0]) begin
          coeffs_719 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_720 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d0 == rs2[9:0]) begin
          coeffs_720 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_721 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d1 == rs2[9:0]) begin
          coeffs_721 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_722 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d2 == rs2[9:0]) begin
          coeffs_722 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_723 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d3 == rs2[9:0]) begin
          coeffs_723 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_724 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d4 == rs2[9:0]) begin
          coeffs_724 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_725 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d5 == rs2[9:0]) begin
          coeffs_725 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_726 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d6 == rs2[9:0]) begin
          coeffs_726 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_727 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d7 == rs2[9:0]) begin
          coeffs_727 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_728 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d8 == rs2[9:0]) begin
          coeffs_728 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_729 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2d9 == rs2[9:0]) begin
          coeffs_729 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_730 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2da == rs2[9:0]) begin
          coeffs_730 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_731 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2db == rs2[9:0]) begin
          coeffs_731 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_732 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2dc == rs2[9:0]) begin
          coeffs_732 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_733 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2dd == rs2[9:0]) begin
          coeffs_733 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_734 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2de == rs2[9:0]) begin
          coeffs_734 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_735 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2df == rs2[9:0]) begin
          coeffs_735 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_736 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e0 == rs2[9:0]) begin
          coeffs_736 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_737 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e1 == rs2[9:0]) begin
          coeffs_737 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_738 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e2 == rs2[9:0]) begin
          coeffs_738 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_739 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e3 == rs2[9:0]) begin
          coeffs_739 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_740 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e4 == rs2[9:0]) begin
          coeffs_740 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_741 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e5 == rs2[9:0]) begin
          coeffs_741 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_742 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e6 == rs2[9:0]) begin
          coeffs_742 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_743 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e7 == rs2[9:0]) begin
          coeffs_743 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_744 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e8 == rs2[9:0]) begin
          coeffs_744 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_745 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2e9 == rs2[9:0]) begin
          coeffs_745 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_746 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ea == rs2[9:0]) begin
          coeffs_746 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_747 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2eb == rs2[9:0]) begin
          coeffs_747 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_748 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ec == rs2[9:0]) begin
          coeffs_748 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_749 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ed == rs2[9:0]) begin
          coeffs_749 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_750 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ee == rs2[9:0]) begin
          coeffs_750 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_751 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ef == rs2[9:0]) begin
          coeffs_751 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_752 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f0 == rs2[9:0]) begin
          coeffs_752 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_753 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f1 == rs2[9:0]) begin
          coeffs_753 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_754 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f2 == rs2[9:0]) begin
          coeffs_754 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_755 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f3 == rs2[9:0]) begin
          coeffs_755 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_756 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f4 == rs2[9:0]) begin
          coeffs_756 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_757 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f5 == rs2[9:0]) begin
          coeffs_757 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_758 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f6 == rs2[9:0]) begin
          coeffs_758 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_759 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f7 == rs2[9:0]) begin
          coeffs_759 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_760 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f8 == rs2[9:0]) begin
          coeffs_760 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_761 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2f9 == rs2[9:0]) begin
          coeffs_761 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_762 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2fa == rs2[9:0]) begin
          coeffs_762 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_763 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2fb == rs2[9:0]) begin
          coeffs_763 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_764 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2fc == rs2[9:0]) begin
          coeffs_764 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_765 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2fd == rs2[9:0]) begin
          coeffs_765 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_766 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2fe == rs2[9:0]) begin
          coeffs_766 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_767 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h2ff == rs2[9:0]) begin
          coeffs_767 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_768 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h300 == rs2[9:0]) begin
          coeffs_768 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_769 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h301 == rs2[9:0]) begin
          coeffs_769 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_770 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h302 == rs2[9:0]) begin
          coeffs_770 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_771 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h303 == rs2[9:0]) begin
          coeffs_771 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_772 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h304 == rs2[9:0]) begin
          coeffs_772 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_773 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h305 == rs2[9:0]) begin
          coeffs_773 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_774 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h306 == rs2[9:0]) begin
          coeffs_774 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_775 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h307 == rs2[9:0]) begin
          coeffs_775 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_776 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h308 == rs2[9:0]) begin
          coeffs_776 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_777 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h309 == rs2[9:0]) begin
          coeffs_777 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_778 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h30a == rs2[9:0]) begin
          coeffs_778 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_779 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h30b == rs2[9:0]) begin
          coeffs_779 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_780 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h30c == rs2[9:0]) begin
          coeffs_780 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_781 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h30d == rs2[9:0]) begin
          coeffs_781 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_782 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h30e == rs2[9:0]) begin
          coeffs_782 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_783 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h30f == rs2[9:0]) begin
          coeffs_783 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_784 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h310 == rs2[9:0]) begin
          coeffs_784 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_785 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h311 == rs2[9:0]) begin
          coeffs_785 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_786 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h312 == rs2[9:0]) begin
          coeffs_786 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_787 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h313 == rs2[9:0]) begin
          coeffs_787 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_788 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h314 == rs2[9:0]) begin
          coeffs_788 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_789 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h315 == rs2[9:0]) begin
          coeffs_789 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_790 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h316 == rs2[9:0]) begin
          coeffs_790 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_791 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h317 == rs2[9:0]) begin
          coeffs_791 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_792 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h318 == rs2[9:0]) begin
          coeffs_792 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_793 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h319 == rs2[9:0]) begin
          coeffs_793 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_794 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h31a == rs2[9:0]) begin
          coeffs_794 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_795 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h31b == rs2[9:0]) begin
          coeffs_795 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_796 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h31c == rs2[9:0]) begin
          coeffs_796 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_797 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h31d == rs2[9:0]) begin
          coeffs_797 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_798 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h31e == rs2[9:0]) begin
          coeffs_798 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_799 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h31f == rs2[9:0]) begin
          coeffs_799 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_800 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h320 == rs2[9:0]) begin
          coeffs_800 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_801 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h321 == rs2[9:0]) begin
          coeffs_801 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_802 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h322 == rs2[9:0]) begin
          coeffs_802 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_803 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h323 == rs2[9:0]) begin
          coeffs_803 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_804 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h324 == rs2[9:0]) begin
          coeffs_804 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_805 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h325 == rs2[9:0]) begin
          coeffs_805 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_806 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h326 == rs2[9:0]) begin
          coeffs_806 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_807 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h327 == rs2[9:0]) begin
          coeffs_807 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_808 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h328 == rs2[9:0]) begin
          coeffs_808 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_809 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h329 == rs2[9:0]) begin
          coeffs_809 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_810 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h32a == rs2[9:0]) begin
          coeffs_810 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_811 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h32b == rs2[9:0]) begin
          coeffs_811 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_812 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h32c == rs2[9:0]) begin
          coeffs_812 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_813 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h32d == rs2[9:0]) begin
          coeffs_813 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_814 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h32e == rs2[9:0]) begin
          coeffs_814 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_815 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h32f == rs2[9:0]) begin
          coeffs_815 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_816 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h330 == rs2[9:0]) begin
          coeffs_816 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_817 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h331 == rs2[9:0]) begin
          coeffs_817 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_818 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h332 == rs2[9:0]) begin
          coeffs_818 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_819 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h333 == rs2[9:0]) begin
          coeffs_819 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_820 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h334 == rs2[9:0]) begin
          coeffs_820 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_821 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h335 == rs2[9:0]) begin
          coeffs_821 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_822 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h336 == rs2[9:0]) begin
          coeffs_822 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_823 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h337 == rs2[9:0]) begin
          coeffs_823 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_824 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h338 == rs2[9:0]) begin
          coeffs_824 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_825 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h339 == rs2[9:0]) begin
          coeffs_825 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_826 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h33a == rs2[9:0]) begin
          coeffs_826 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_827 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h33b == rs2[9:0]) begin
          coeffs_827 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_828 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h33c == rs2[9:0]) begin
          coeffs_828 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_829 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h33d == rs2[9:0]) begin
          coeffs_829 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_830 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h33e == rs2[9:0]) begin
          coeffs_830 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_831 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h33f == rs2[9:0]) begin
          coeffs_831 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_832 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h340 == rs2[9:0]) begin
          coeffs_832 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_833 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h341 == rs2[9:0]) begin
          coeffs_833 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_834 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h342 == rs2[9:0]) begin
          coeffs_834 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_835 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h343 == rs2[9:0]) begin
          coeffs_835 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_836 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h344 == rs2[9:0]) begin
          coeffs_836 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_837 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h345 == rs2[9:0]) begin
          coeffs_837 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_838 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h346 == rs2[9:0]) begin
          coeffs_838 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_839 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h347 == rs2[9:0]) begin
          coeffs_839 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_840 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h348 == rs2[9:0]) begin
          coeffs_840 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_841 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h349 == rs2[9:0]) begin
          coeffs_841 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_842 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h34a == rs2[9:0]) begin
          coeffs_842 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_843 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h34b == rs2[9:0]) begin
          coeffs_843 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_844 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h34c == rs2[9:0]) begin
          coeffs_844 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_845 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h34d == rs2[9:0]) begin
          coeffs_845 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_846 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h34e == rs2[9:0]) begin
          coeffs_846 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_847 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h34f == rs2[9:0]) begin
          coeffs_847 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_848 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h350 == rs2[9:0]) begin
          coeffs_848 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_849 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h351 == rs2[9:0]) begin
          coeffs_849 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_850 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h352 == rs2[9:0]) begin
          coeffs_850 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_851 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h353 == rs2[9:0]) begin
          coeffs_851 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_852 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h354 == rs2[9:0]) begin
          coeffs_852 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_853 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h355 == rs2[9:0]) begin
          coeffs_853 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_854 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h356 == rs2[9:0]) begin
          coeffs_854 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_855 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h357 == rs2[9:0]) begin
          coeffs_855 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_856 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h358 == rs2[9:0]) begin
          coeffs_856 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_857 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h359 == rs2[9:0]) begin
          coeffs_857 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_858 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h35a == rs2[9:0]) begin
          coeffs_858 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_859 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h35b == rs2[9:0]) begin
          coeffs_859 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_860 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h35c == rs2[9:0]) begin
          coeffs_860 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_861 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h35d == rs2[9:0]) begin
          coeffs_861 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_862 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h35e == rs2[9:0]) begin
          coeffs_862 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_863 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h35f == rs2[9:0]) begin
          coeffs_863 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_864 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h360 == rs2[9:0]) begin
          coeffs_864 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_865 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h361 == rs2[9:0]) begin
          coeffs_865 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_866 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h362 == rs2[9:0]) begin
          coeffs_866 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_867 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h363 == rs2[9:0]) begin
          coeffs_867 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_868 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h364 == rs2[9:0]) begin
          coeffs_868 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_869 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h365 == rs2[9:0]) begin
          coeffs_869 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_870 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h366 == rs2[9:0]) begin
          coeffs_870 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_871 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h367 == rs2[9:0]) begin
          coeffs_871 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_872 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h368 == rs2[9:0]) begin
          coeffs_872 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_873 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h369 == rs2[9:0]) begin
          coeffs_873 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_874 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h36a == rs2[9:0]) begin
          coeffs_874 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_875 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h36b == rs2[9:0]) begin
          coeffs_875 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_876 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h36c == rs2[9:0]) begin
          coeffs_876 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_877 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h36d == rs2[9:0]) begin
          coeffs_877 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_878 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h36e == rs2[9:0]) begin
          coeffs_878 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_879 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h36f == rs2[9:0]) begin
          coeffs_879 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_880 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h370 == rs2[9:0]) begin
          coeffs_880 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_881 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h371 == rs2[9:0]) begin
          coeffs_881 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_882 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h372 == rs2[9:0]) begin
          coeffs_882 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_883 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h373 == rs2[9:0]) begin
          coeffs_883 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_884 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h374 == rs2[9:0]) begin
          coeffs_884 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_885 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h375 == rs2[9:0]) begin
          coeffs_885 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_886 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h376 == rs2[9:0]) begin
          coeffs_886 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_887 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h377 == rs2[9:0]) begin
          coeffs_887 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_888 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h378 == rs2[9:0]) begin
          coeffs_888 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_889 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h379 == rs2[9:0]) begin
          coeffs_889 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_890 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h37a == rs2[9:0]) begin
          coeffs_890 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_891 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h37b == rs2[9:0]) begin
          coeffs_891 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_892 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h37c == rs2[9:0]) begin
          coeffs_892 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_893 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h37d == rs2[9:0]) begin
          coeffs_893 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_894 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h37e == rs2[9:0]) begin
          coeffs_894 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_895 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h37f == rs2[9:0]) begin
          coeffs_895 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_896 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h380 == rs2[9:0]) begin
          coeffs_896 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_897 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h381 == rs2[9:0]) begin
          coeffs_897 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_898 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h382 == rs2[9:0]) begin
          coeffs_898 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_899 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h383 == rs2[9:0]) begin
          coeffs_899 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_900 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h384 == rs2[9:0]) begin
          coeffs_900 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_901 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h385 == rs2[9:0]) begin
          coeffs_901 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_902 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h386 == rs2[9:0]) begin
          coeffs_902 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_903 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h387 == rs2[9:0]) begin
          coeffs_903 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_904 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h388 == rs2[9:0]) begin
          coeffs_904 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_905 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h389 == rs2[9:0]) begin
          coeffs_905 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_906 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h38a == rs2[9:0]) begin
          coeffs_906 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_907 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h38b == rs2[9:0]) begin
          coeffs_907 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_908 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h38c == rs2[9:0]) begin
          coeffs_908 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_909 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h38d == rs2[9:0]) begin
          coeffs_909 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_910 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h38e == rs2[9:0]) begin
          coeffs_910 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_911 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h38f == rs2[9:0]) begin
          coeffs_911 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_912 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h390 == rs2[9:0]) begin
          coeffs_912 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_913 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h391 == rs2[9:0]) begin
          coeffs_913 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_914 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h392 == rs2[9:0]) begin
          coeffs_914 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_915 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h393 == rs2[9:0]) begin
          coeffs_915 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_916 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h394 == rs2[9:0]) begin
          coeffs_916 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_917 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h395 == rs2[9:0]) begin
          coeffs_917 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_918 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h396 == rs2[9:0]) begin
          coeffs_918 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_919 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h397 == rs2[9:0]) begin
          coeffs_919 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_920 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h398 == rs2[9:0]) begin
          coeffs_920 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_921 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h399 == rs2[9:0]) begin
          coeffs_921 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_922 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h39a == rs2[9:0]) begin
          coeffs_922 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_923 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h39b == rs2[9:0]) begin
          coeffs_923 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_924 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h39c == rs2[9:0]) begin
          coeffs_924 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_925 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h39d == rs2[9:0]) begin
          coeffs_925 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_926 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h39e == rs2[9:0]) begin
          coeffs_926 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_927 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h39f == rs2[9:0]) begin
          coeffs_927 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_928 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a0 == rs2[9:0]) begin
          coeffs_928 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_929 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a1 == rs2[9:0]) begin
          coeffs_929 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_930 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a2 == rs2[9:0]) begin
          coeffs_930 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_931 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a3 == rs2[9:0]) begin
          coeffs_931 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_932 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a4 == rs2[9:0]) begin
          coeffs_932 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_933 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a5 == rs2[9:0]) begin
          coeffs_933 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_934 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a6 == rs2[9:0]) begin
          coeffs_934 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_935 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a7 == rs2[9:0]) begin
          coeffs_935 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_936 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a8 == rs2[9:0]) begin
          coeffs_936 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_937 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3a9 == rs2[9:0]) begin
          coeffs_937 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_938 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3aa == rs2[9:0]) begin
          coeffs_938 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_939 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3ab == rs2[9:0]) begin
          coeffs_939 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_940 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3ac == rs2[9:0]) begin
          coeffs_940 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_941 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3ad == rs2[9:0]) begin
          coeffs_941 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_942 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3ae == rs2[9:0]) begin
          coeffs_942 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_943 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3af == rs2[9:0]) begin
          coeffs_943 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_944 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b0 == rs2[9:0]) begin
          coeffs_944 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_945 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b1 == rs2[9:0]) begin
          coeffs_945 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_946 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b2 == rs2[9:0]) begin
          coeffs_946 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_947 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b3 == rs2[9:0]) begin
          coeffs_947 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_948 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b4 == rs2[9:0]) begin
          coeffs_948 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_949 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b5 == rs2[9:0]) begin
          coeffs_949 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_950 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b6 == rs2[9:0]) begin
          coeffs_950 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_951 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b7 == rs2[9:0]) begin
          coeffs_951 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_952 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b8 == rs2[9:0]) begin
          coeffs_952 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_953 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3b9 == rs2[9:0]) begin
          coeffs_953 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_954 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3ba == rs2[9:0]) begin
          coeffs_954 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_955 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3bb == rs2[9:0]) begin
          coeffs_955 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_956 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3bc == rs2[9:0]) begin
          coeffs_956 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_957 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3bd == rs2[9:0]) begin
          coeffs_957 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_958 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3be == rs2[9:0]) begin
          coeffs_958 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_959 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3bf == rs2[9:0]) begin
          coeffs_959 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_960 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c0 == rs2[9:0]) begin
          coeffs_960 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_961 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c1 == rs2[9:0]) begin
          coeffs_961 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_962 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c2 == rs2[9:0]) begin
          coeffs_962 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_963 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c3 == rs2[9:0]) begin
          coeffs_963 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_964 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c4 == rs2[9:0]) begin
          coeffs_964 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_965 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c5 == rs2[9:0]) begin
          coeffs_965 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_966 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c6 == rs2[9:0]) begin
          coeffs_966 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_967 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c7 == rs2[9:0]) begin
          coeffs_967 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_968 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c8 == rs2[9:0]) begin
          coeffs_968 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_969 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3c9 == rs2[9:0]) begin
          coeffs_969 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_970 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3ca == rs2[9:0]) begin
          coeffs_970 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_971 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3cb == rs2[9:0]) begin
          coeffs_971 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_972 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3cc == rs2[9:0]) begin
          coeffs_972 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_973 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3cd == rs2[9:0]) begin
          coeffs_973 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_974 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3ce == rs2[9:0]) begin
          coeffs_974 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_975 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3cf == rs2[9:0]) begin
          coeffs_975 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_976 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d0 == rs2[9:0]) begin
          coeffs_976 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_977 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d1 == rs2[9:0]) begin
          coeffs_977 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_978 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d2 == rs2[9:0]) begin
          coeffs_978 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_979 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d3 == rs2[9:0]) begin
          coeffs_979 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_980 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d4 == rs2[9:0]) begin
          coeffs_980 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_981 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d5 == rs2[9:0]) begin
          coeffs_981 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_982 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d6 == rs2[9:0]) begin
          coeffs_982 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_983 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d7 == rs2[9:0]) begin
          coeffs_983 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_984 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d8 == rs2[9:0]) begin
          coeffs_984 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_985 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3d9 == rs2[9:0]) begin
          coeffs_985 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_986 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3da == rs2[9:0]) begin
          coeffs_986 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_987 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3db == rs2[9:0]) begin
          coeffs_987 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_988 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3dc == rs2[9:0]) begin
          coeffs_988 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_989 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3dd == rs2[9:0]) begin
          coeffs_989 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_990 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3de == rs2[9:0]) begin
          coeffs_990 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_991 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3df == rs2[9:0]) begin
          coeffs_991 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_992 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3e0 == rs2[9:0]) begin
          coeffs_992 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_993 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3e1 == rs2[9:0]) begin
          coeffs_993 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_994 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3e2 == rs2[9:0]) begin
          coeffs_994 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_995 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3e3 == rs2[9:0]) begin
          coeffs_995 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_996 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3e4 == rs2[9:0]) begin
          coeffs_996 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_997 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3e5 == rs2[9:0]) begin
          coeffs_997 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_998 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3e6 == rs2[9:0]) begin
          coeffs_998 <= rs1;
        end
      end
    end
    if (reset) begin
      coeffs_999 <= 32'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        if (10'h3e7 == rs2[9:0]) begin
          coeffs_999 <= rs1;
        end
      end
    end
    if (reset) begin
      data_0 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_0 <= rs1;
        end
      end
    end
    if (reset) begin
      data_1 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_1 <= data_0;
        end
      end
    end
    if (reset) begin
      data_2 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_2 <= data_1;
        end
      end
    end
    if (reset) begin
      data_3 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_3 <= data_2;
        end
      end
    end
    if (reset) begin
      data_4 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_4 <= data_3;
        end
      end
    end
    if (reset) begin
      data_5 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_5 <= data_4;
        end
      end
    end
    if (reset) begin
      data_6 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_6 <= data_5;
        end
      end
    end
    if (reset) begin
      data_7 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_7 <= data_6;
        end
      end
    end
    if (reset) begin
      data_8 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_8 <= data_7;
        end
      end
    end
    if (reset) begin
      data_9 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_9 <= data_8;
        end
      end
    end
    if (reset) begin
      data_10 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_10 <= data_9;
        end
      end
    end
    if (reset) begin
      data_11 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_11 <= data_10;
        end
      end
    end
    if (reset) begin
      data_12 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_12 <= data_11;
        end
      end
    end
    if (reset) begin
      data_13 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_13 <= data_12;
        end
      end
    end
    if (reset) begin
      data_14 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_14 <= data_13;
        end
      end
    end
    if (reset) begin
      data_15 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_15 <= data_14;
        end
      end
    end
    if (reset) begin
      data_16 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_16 <= data_15;
        end
      end
    end
    if (reset) begin
      data_17 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_17 <= data_16;
        end
      end
    end
    if (reset) begin
      data_18 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_18 <= data_17;
        end
      end
    end
    if (reset) begin
      data_19 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_19 <= data_18;
        end
      end
    end
    if (reset) begin
      data_20 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_20 <= data_19;
        end
      end
    end
    if (reset) begin
      data_21 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_21 <= data_20;
        end
      end
    end
    if (reset) begin
      data_22 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_22 <= data_21;
        end
      end
    end
    if (reset) begin
      data_23 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_23 <= data_22;
        end
      end
    end
    if (reset) begin
      data_24 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_24 <= data_23;
        end
      end
    end
    if (reset) begin
      data_25 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_25 <= data_24;
        end
      end
    end
    if (reset) begin
      data_26 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_26 <= data_25;
        end
      end
    end
    if (reset) begin
      data_27 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_27 <= data_26;
        end
      end
    end
    if (reset) begin
      data_28 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_28 <= data_27;
        end
      end
    end
    if (reset) begin
      data_29 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_29 <= data_28;
        end
      end
    end
    if (reset) begin
      data_30 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_30 <= data_29;
        end
      end
    end
    if (reset) begin
      data_31 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_31 <= data_30;
        end
      end
    end
    if (reset) begin
      data_32 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_32 <= data_31;
        end
      end
    end
    if (reset) begin
      data_33 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_33 <= data_32;
        end
      end
    end
    if (reset) begin
      data_34 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_34 <= data_33;
        end
      end
    end
    if (reset) begin
      data_35 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_35 <= data_34;
        end
      end
    end
    if (reset) begin
      data_36 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_36 <= data_35;
        end
      end
    end
    if (reset) begin
      data_37 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_37 <= data_36;
        end
      end
    end
    if (reset) begin
      data_38 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_38 <= data_37;
        end
      end
    end
    if (reset) begin
      data_39 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_39 <= data_38;
        end
      end
    end
    if (reset) begin
      data_40 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_40 <= data_39;
        end
      end
    end
    if (reset) begin
      data_41 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_41 <= data_40;
        end
      end
    end
    if (reset) begin
      data_42 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_42 <= data_41;
        end
      end
    end
    if (reset) begin
      data_43 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_43 <= data_42;
        end
      end
    end
    if (reset) begin
      data_44 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_44 <= data_43;
        end
      end
    end
    if (reset) begin
      data_45 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_45 <= data_44;
        end
      end
    end
    if (reset) begin
      data_46 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_46 <= data_45;
        end
      end
    end
    if (reset) begin
      data_47 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_47 <= data_46;
        end
      end
    end
    if (reset) begin
      data_48 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_48 <= data_47;
        end
      end
    end
    if (reset) begin
      data_49 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_49 <= data_48;
        end
      end
    end
    if (reset) begin
      data_50 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_50 <= data_49;
        end
      end
    end
    if (reset) begin
      data_51 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_51 <= data_50;
        end
      end
    end
    if (reset) begin
      data_52 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_52 <= data_51;
        end
      end
    end
    if (reset) begin
      data_53 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_53 <= data_52;
        end
      end
    end
    if (reset) begin
      data_54 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_54 <= data_53;
        end
      end
    end
    if (reset) begin
      data_55 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_55 <= data_54;
        end
      end
    end
    if (reset) begin
      data_56 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_56 <= data_55;
        end
      end
    end
    if (reset) begin
      data_57 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_57 <= data_56;
        end
      end
    end
    if (reset) begin
      data_58 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_58 <= data_57;
        end
      end
    end
    if (reset) begin
      data_59 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_59 <= data_58;
        end
      end
    end
    if (reset) begin
      data_60 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_60 <= data_59;
        end
      end
    end
    if (reset) begin
      data_61 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_61 <= data_60;
        end
      end
    end
    if (reset) begin
      data_62 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_62 <= data_61;
        end
      end
    end
    if (reset) begin
      data_63 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_63 <= data_62;
        end
      end
    end
    if (reset) begin
      data_64 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_64 <= data_63;
        end
      end
    end
    if (reset) begin
      data_65 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_65 <= data_64;
        end
      end
    end
    if (reset) begin
      data_66 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_66 <= data_65;
        end
      end
    end
    if (reset) begin
      data_67 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_67 <= data_66;
        end
      end
    end
    if (reset) begin
      data_68 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_68 <= data_67;
        end
      end
    end
    if (reset) begin
      data_69 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_69 <= data_68;
        end
      end
    end
    if (reset) begin
      data_70 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_70 <= data_69;
        end
      end
    end
    if (reset) begin
      data_71 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_71 <= data_70;
        end
      end
    end
    if (reset) begin
      data_72 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_72 <= data_71;
        end
      end
    end
    if (reset) begin
      data_73 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_73 <= data_72;
        end
      end
    end
    if (reset) begin
      data_74 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_74 <= data_73;
        end
      end
    end
    if (reset) begin
      data_75 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_75 <= data_74;
        end
      end
    end
    if (reset) begin
      data_76 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_76 <= data_75;
        end
      end
    end
    if (reset) begin
      data_77 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_77 <= data_76;
        end
      end
    end
    if (reset) begin
      data_78 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_78 <= data_77;
        end
      end
    end
    if (reset) begin
      data_79 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_79 <= data_78;
        end
      end
    end
    if (reset) begin
      data_80 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_80 <= data_79;
        end
      end
    end
    if (reset) begin
      data_81 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_81 <= data_80;
        end
      end
    end
    if (reset) begin
      data_82 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_82 <= data_81;
        end
      end
    end
    if (reset) begin
      data_83 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_83 <= data_82;
        end
      end
    end
    if (reset) begin
      data_84 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_84 <= data_83;
        end
      end
    end
    if (reset) begin
      data_85 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_85 <= data_84;
        end
      end
    end
    if (reset) begin
      data_86 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_86 <= data_85;
        end
      end
    end
    if (reset) begin
      data_87 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_87 <= data_86;
        end
      end
    end
    if (reset) begin
      data_88 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_88 <= data_87;
        end
      end
    end
    if (reset) begin
      data_89 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_89 <= data_88;
        end
      end
    end
    if (reset) begin
      data_90 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_90 <= data_89;
        end
      end
    end
    if (reset) begin
      data_91 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_91 <= data_90;
        end
      end
    end
    if (reset) begin
      data_92 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_92 <= data_91;
        end
      end
    end
    if (reset) begin
      data_93 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_93 <= data_92;
        end
      end
    end
    if (reset) begin
      data_94 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_94 <= data_93;
        end
      end
    end
    if (reset) begin
      data_95 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_95 <= data_94;
        end
      end
    end
    if (reset) begin
      data_96 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_96 <= data_95;
        end
      end
    end
    if (reset) begin
      data_97 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_97 <= data_96;
        end
      end
    end
    if (reset) begin
      data_98 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_98 <= data_97;
        end
      end
    end
    if (reset) begin
      data_99 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_99 <= data_98;
        end
      end
    end
    if (reset) begin
      data_100 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_100 <= data_99;
        end
      end
    end
    if (reset) begin
      data_101 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_101 <= data_100;
        end
      end
    end
    if (reset) begin
      data_102 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_102 <= data_101;
        end
      end
    end
    if (reset) begin
      data_103 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_103 <= data_102;
        end
      end
    end
    if (reset) begin
      data_104 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_104 <= data_103;
        end
      end
    end
    if (reset) begin
      data_105 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_105 <= data_104;
        end
      end
    end
    if (reset) begin
      data_106 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_106 <= data_105;
        end
      end
    end
    if (reset) begin
      data_107 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_107 <= data_106;
        end
      end
    end
    if (reset) begin
      data_108 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_108 <= data_107;
        end
      end
    end
    if (reset) begin
      data_109 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_109 <= data_108;
        end
      end
    end
    if (reset) begin
      data_110 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_110 <= data_109;
        end
      end
    end
    if (reset) begin
      data_111 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_111 <= data_110;
        end
      end
    end
    if (reset) begin
      data_112 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_112 <= data_111;
        end
      end
    end
    if (reset) begin
      data_113 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_113 <= data_112;
        end
      end
    end
    if (reset) begin
      data_114 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_114 <= data_113;
        end
      end
    end
    if (reset) begin
      data_115 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_115 <= data_114;
        end
      end
    end
    if (reset) begin
      data_116 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_116 <= data_115;
        end
      end
    end
    if (reset) begin
      data_117 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_117 <= data_116;
        end
      end
    end
    if (reset) begin
      data_118 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_118 <= data_117;
        end
      end
    end
    if (reset) begin
      data_119 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_119 <= data_118;
        end
      end
    end
    if (reset) begin
      data_120 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_120 <= data_119;
        end
      end
    end
    if (reset) begin
      data_121 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_121 <= data_120;
        end
      end
    end
    if (reset) begin
      data_122 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_122 <= data_121;
        end
      end
    end
    if (reset) begin
      data_123 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_123 <= data_122;
        end
      end
    end
    if (reset) begin
      data_124 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_124 <= data_123;
        end
      end
    end
    if (reset) begin
      data_125 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_125 <= data_124;
        end
      end
    end
    if (reset) begin
      data_126 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_126 <= data_125;
        end
      end
    end
    if (reset) begin
      data_127 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_127 <= data_126;
        end
      end
    end
    if (reset) begin
      data_128 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_128 <= data_127;
        end
      end
    end
    if (reset) begin
      data_129 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_129 <= data_128;
        end
      end
    end
    if (reset) begin
      data_130 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_130 <= data_129;
        end
      end
    end
    if (reset) begin
      data_131 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_131 <= data_130;
        end
      end
    end
    if (reset) begin
      data_132 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_132 <= data_131;
        end
      end
    end
    if (reset) begin
      data_133 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_133 <= data_132;
        end
      end
    end
    if (reset) begin
      data_134 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_134 <= data_133;
        end
      end
    end
    if (reset) begin
      data_135 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_135 <= data_134;
        end
      end
    end
    if (reset) begin
      data_136 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_136 <= data_135;
        end
      end
    end
    if (reset) begin
      data_137 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_137 <= data_136;
        end
      end
    end
    if (reset) begin
      data_138 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_138 <= data_137;
        end
      end
    end
    if (reset) begin
      data_139 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_139 <= data_138;
        end
      end
    end
    if (reset) begin
      data_140 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_140 <= data_139;
        end
      end
    end
    if (reset) begin
      data_141 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_141 <= data_140;
        end
      end
    end
    if (reset) begin
      data_142 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_142 <= data_141;
        end
      end
    end
    if (reset) begin
      data_143 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_143 <= data_142;
        end
      end
    end
    if (reset) begin
      data_144 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_144 <= data_143;
        end
      end
    end
    if (reset) begin
      data_145 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_145 <= data_144;
        end
      end
    end
    if (reset) begin
      data_146 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_146 <= data_145;
        end
      end
    end
    if (reset) begin
      data_147 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_147 <= data_146;
        end
      end
    end
    if (reset) begin
      data_148 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_148 <= data_147;
        end
      end
    end
    if (reset) begin
      data_149 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_149 <= data_148;
        end
      end
    end
    if (reset) begin
      data_150 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_150 <= data_149;
        end
      end
    end
    if (reset) begin
      data_151 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_151 <= data_150;
        end
      end
    end
    if (reset) begin
      data_152 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_152 <= data_151;
        end
      end
    end
    if (reset) begin
      data_153 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_153 <= data_152;
        end
      end
    end
    if (reset) begin
      data_154 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_154 <= data_153;
        end
      end
    end
    if (reset) begin
      data_155 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_155 <= data_154;
        end
      end
    end
    if (reset) begin
      data_156 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_156 <= data_155;
        end
      end
    end
    if (reset) begin
      data_157 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_157 <= data_156;
        end
      end
    end
    if (reset) begin
      data_158 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_158 <= data_157;
        end
      end
    end
    if (reset) begin
      data_159 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_159 <= data_158;
        end
      end
    end
    if (reset) begin
      data_160 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_160 <= data_159;
        end
      end
    end
    if (reset) begin
      data_161 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_161 <= data_160;
        end
      end
    end
    if (reset) begin
      data_162 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_162 <= data_161;
        end
      end
    end
    if (reset) begin
      data_163 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_163 <= data_162;
        end
      end
    end
    if (reset) begin
      data_164 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_164 <= data_163;
        end
      end
    end
    if (reset) begin
      data_165 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_165 <= data_164;
        end
      end
    end
    if (reset) begin
      data_166 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_166 <= data_165;
        end
      end
    end
    if (reset) begin
      data_167 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_167 <= data_166;
        end
      end
    end
    if (reset) begin
      data_168 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_168 <= data_167;
        end
      end
    end
    if (reset) begin
      data_169 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_169 <= data_168;
        end
      end
    end
    if (reset) begin
      data_170 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_170 <= data_169;
        end
      end
    end
    if (reset) begin
      data_171 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_171 <= data_170;
        end
      end
    end
    if (reset) begin
      data_172 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_172 <= data_171;
        end
      end
    end
    if (reset) begin
      data_173 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_173 <= data_172;
        end
      end
    end
    if (reset) begin
      data_174 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_174 <= data_173;
        end
      end
    end
    if (reset) begin
      data_175 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_175 <= data_174;
        end
      end
    end
    if (reset) begin
      data_176 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_176 <= data_175;
        end
      end
    end
    if (reset) begin
      data_177 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_177 <= data_176;
        end
      end
    end
    if (reset) begin
      data_178 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_178 <= data_177;
        end
      end
    end
    if (reset) begin
      data_179 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_179 <= data_178;
        end
      end
    end
    if (reset) begin
      data_180 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_180 <= data_179;
        end
      end
    end
    if (reset) begin
      data_181 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_181 <= data_180;
        end
      end
    end
    if (reset) begin
      data_182 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_182 <= data_181;
        end
      end
    end
    if (reset) begin
      data_183 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_183 <= data_182;
        end
      end
    end
    if (reset) begin
      data_184 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_184 <= data_183;
        end
      end
    end
    if (reset) begin
      data_185 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_185 <= data_184;
        end
      end
    end
    if (reset) begin
      data_186 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_186 <= data_185;
        end
      end
    end
    if (reset) begin
      data_187 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_187 <= data_186;
        end
      end
    end
    if (reset) begin
      data_188 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_188 <= data_187;
        end
      end
    end
    if (reset) begin
      data_189 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_189 <= data_188;
        end
      end
    end
    if (reset) begin
      data_190 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_190 <= data_189;
        end
      end
    end
    if (reset) begin
      data_191 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_191 <= data_190;
        end
      end
    end
    if (reset) begin
      data_192 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_192 <= data_191;
        end
      end
    end
    if (reset) begin
      data_193 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_193 <= data_192;
        end
      end
    end
    if (reset) begin
      data_194 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_194 <= data_193;
        end
      end
    end
    if (reset) begin
      data_195 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_195 <= data_194;
        end
      end
    end
    if (reset) begin
      data_196 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_196 <= data_195;
        end
      end
    end
    if (reset) begin
      data_197 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_197 <= data_196;
        end
      end
    end
    if (reset) begin
      data_198 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_198 <= data_197;
        end
      end
    end
    if (reset) begin
      data_199 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_199 <= data_198;
        end
      end
    end
    if (reset) begin
      data_200 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_200 <= data_199;
        end
      end
    end
    if (reset) begin
      data_201 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_201 <= data_200;
        end
      end
    end
    if (reset) begin
      data_202 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_202 <= data_201;
        end
      end
    end
    if (reset) begin
      data_203 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_203 <= data_202;
        end
      end
    end
    if (reset) begin
      data_204 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_204 <= data_203;
        end
      end
    end
    if (reset) begin
      data_205 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_205 <= data_204;
        end
      end
    end
    if (reset) begin
      data_206 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_206 <= data_205;
        end
      end
    end
    if (reset) begin
      data_207 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_207 <= data_206;
        end
      end
    end
    if (reset) begin
      data_208 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_208 <= data_207;
        end
      end
    end
    if (reset) begin
      data_209 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_209 <= data_208;
        end
      end
    end
    if (reset) begin
      data_210 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_210 <= data_209;
        end
      end
    end
    if (reset) begin
      data_211 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_211 <= data_210;
        end
      end
    end
    if (reset) begin
      data_212 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_212 <= data_211;
        end
      end
    end
    if (reset) begin
      data_213 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_213 <= data_212;
        end
      end
    end
    if (reset) begin
      data_214 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_214 <= data_213;
        end
      end
    end
    if (reset) begin
      data_215 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_215 <= data_214;
        end
      end
    end
    if (reset) begin
      data_216 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_216 <= data_215;
        end
      end
    end
    if (reset) begin
      data_217 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_217 <= data_216;
        end
      end
    end
    if (reset) begin
      data_218 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_218 <= data_217;
        end
      end
    end
    if (reset) begin
      data_219 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_219 <= data_218;
        end
      end
    end
    if (reset) begin
      data_220 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_220 <= data_219;
        end
      end
    end
    if (reset) begin
      data_221 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_221 <= data_220;
        end
      end
    end
    if (reset) begin
      data_222 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_222 <= data_221;
        end
      end
    end
    if (reset) begin
      data_223 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_223 <= data_222;
        end
      end
    end
    if (reset) begin
      data_224 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_224 <= data_223;
        end
      end
    end
    if (reset) begin
      data_225 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_225 <= data_224;
        end
      end
    end
    if (reset) begin
      data_226 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_226 <= data_225;
        end
      end
    end
    if (reset) begin
      data_227 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_227 <= data_226;
        end
      end
    end
    if (reset) begin
      data_228 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_228 <= data_227;
        end
      end
    end
    if (reset) begin
      data_229 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_229 <= data_228;
        end
      end
    end
    if (reset) begin
      data_230 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_230 <= data_229;
        end
      end
    end
    if (reset) begin
      data_231 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_231 <= data_230;
        end
      end
    end
    if (reset) begin
      data_232 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_232 <= data_231;
        end
      end
    end
    if (reset) begin
      data_233 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_233 <= data_232;
        end
      end
    end
    if (reset) begin
      data_234 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_234 <= data_233;
        end
      end
    end
    if (reset) begin
      data_235 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_235 <= data_234;
        end
      end
    end
    if (reset) begin
      data_236 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_236 <= data_235;
        end
      end
    end
    if (reset) begin
      data_237 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_237 <= data_236;
        end
      end
    end
    if (reset) begin
      data_238 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_238 <= data_237;
        end
      end
    end
    if (reset) begin
      data_239 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_239 <= data_238;
        end
      end
    end
    if (reset) begin
      data_240 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_240 <= data_239;
        end
      end
    end
    if (reset) begin
      data_241 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_241 <= data_240;
        end
      end
    end
    if (reset) begin
      data_242 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_242 <= data_241;
        end
      end
    end
    if (reset) begin
      data_243 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_243 <= data_242;
        end
      end
    end
    if (reset) begin
      data_244 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_244 <= data_243;
        end
      end
    end
    if (reset) begin
      data_245 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_245 <= data_244;
        end
      end
    end
    if (reset) begin
      data_246 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_246 <= data_245;
        end
      end
    end
    if (reset) begin
      data_247 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_247 <= data_246;
        end
      end
    end
    if (reset) begin
      data_248 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_248 <= data_247;
        end
      end
    end
    if (reset) begin
      data_249 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_249 <= data_248;
        end
      end
    end
    if (reset) begin
      data_250 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_250 <= data_249;
        end
      end
    end
    if (reset) begin
      data_251 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_251 <= data_250;
        end
      end
    end
    if (reset) begin
      data_252 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_252 <= data_251;
        end
      end
    end
    if (reset) begin
      data_253 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_253 <= data_252;
        end
      end
    end
    if (reset) begin
      data_254 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_254 <= data_253;
        end
      end
    end
    if (reset) begin
      data_255 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_255 <= data_254;
        end
      end
    end
    if (reset) begin
      data_256 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_256 <= data_255;
        end
      end
    end
    if (reset) begin
      data_257 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_257 <= data_256;
        end
      end
    end
    if (reset) begin
      data_258 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_258 <= data_257;
        end
      end
    end
    if (reset) begin
      data_259 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_259 <= data_258;
        end
      end
    end
    if (reset) begin
      data_260 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_260 <= data_259;
        end
      end
    end
    if (reset) begin
      data_261 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_261 <= data_260;
        end
      end
    end
    if (reset) begin
      data_262 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_262 <= data_261;
        end
      end
    end
    if (reset) begin
      data_263 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_263 <= data_262;
        end
      end
    end
    if (reset) begin
      data_264 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_264 <= data_263;
        end
      end
    end
    if (reset) begin
      data_265 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_265 <= data_264;
        end
      end
    end
    if (reset) begin
      data_266 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_266 <= data_265;
        end
      end
    end
    if (reset) begin
      data_267 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_267 <= data_266;
        end
      end
    end
    if (reset) begin
      data_268 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_268 <= data_267;
        end
      end
    end
    if (reset) begin
      data_269 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_269 <= data_268;
        end
      end
    end
    if (reset) begin
      data_270 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_270 <= data_269;
        end
      end
    end
    if (reset) begin
      data_271 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_271 <= data_270;
        end
      end
    end
    if (reset) begin
      data_272 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_272 <= data_271;
        end
      end
    end
    if (reset) begin
      data_273 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_273 <= data_272;
        end
      end
    end
    if (reset) begin
      data_274 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_274 <= data_273;
        end
      end
    end
    if (reset) begin
      data_275 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_275 <= data_274;
        end
      end
    end
    if (reset) begin
      data_276 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_276 <= data_275;
        end
      end
    end
    if (reset) begin
      data_277 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_277 <= data_276;
        end
      end
    end
    if (reset) begin
      data_278 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_278 <= data_277;
        end
      end
    end
    if (reset) begin
      data_279 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_279 <= data_278;
        end
      end
    end
    if (reset) begin
      data_280 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_280 <= data_279;
        end
      end
    end
    if (reset) begin
      data_281 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_281 <= data_280;
        end
      end
    end
    if (reset) begin
      data_282 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_282 <= data_281;
        end
      end
    end
    if (reset) begin
      data_283 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_283 <= data_282;
        end
      end
    end
    if (reset) begin
      data_284 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_284 <= data_283;
        end
      end
    end
    if (reset) begin
      data_285 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_285 <= data_284;
        end
      end
    end
    if (reset) begin
      data_286 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_286 <= data_285;
        end
      end
    end
    if (reset) begin
      data_287 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_287 <= data_286;
        end
      end
    end
    if (reset) begin
      data_288 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_288 <= data_287;
        end
      end
    end
    if (reset) begin
      data_289 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_289 <= data_288;
        end
      end
    end
    if (reset) begin
      data_290 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_290 <= data_289;
        end
      end
    end
    if (reset) begin
      data_291 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_291 <= data_290;
        end
      end
    end
    if (reset) begin
      data_292 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_292 <= data_291;
        end
      end
    end
    if (reset) begin
      data_293 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_293 <= data_292;
        end
      end
    end
    if (reset) begin
      data_294 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_294 <= data_293;
        end
      end
    end
    if (reset) begin
      data_295 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_295 <= data_294;
        end
      end
    end
    if (reset) begin
      data_296 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_296 <= data_295;
        end
      end
    end
    if (reset) begin
      data_297 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_297 <= data_296;
        end
      end
    end
    if (reset) begin
      data_298 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_298 <= data_297;
        end
      end
    end
    if (reset) begin
      data_299 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_299 <= data_298;
        end
      end
    end
    if (reset) begin
      data_300 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_300 <= data_299;
        end
      end
    end
    if (reset) begin
      data_301 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_301 <= data_300;
        end
      end
    end
    if (reset) begin
      data_302 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_302 <= data_301;
        end
      end
    end
    if (reset) begin
      data_303 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_303 <= data_302;
        end
      end
    end
    if (reset) begin
      data_304 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_304 <= data_303;
        end
      end
    end
    if (reset) begin
      data_305 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_305 <= data_304;
        end
      end
    end
    if (reset) begin
      data_306 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_306 <= data_305;
        end
      end
    end
    if (reset) begin
      data_307 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_307 <= data_306;
        end
      end
    end
    if (reset) begin
      data_308 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_308 <= data_307;
        end
      end
    end
    if (reset) begin
      data_309 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_309 <= data_308;
        end
      end
    end
    if (reset) begin
      data_310 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_310 <= data_309;
        end
      end
    end
    if (reset) begin
      data_311 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_311 <= data_310;
        end
      end
    end
    if (reset) begin
      data_312 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_312 <= data_311;
        end
      end
    end
    if (reset) begin
      data_313 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_313 <= data_312;
        end
      end
    end
    if (reset) begin
      data_314 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_314 <= data_313;
        end
      end
    end
    if (reset) begin
      data_315 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_315 <= data_314;
        end
      end
    end
    if (reset) begin
      data_316 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_316 <= data_315;
        end
      end
    end
    if (reset) begin
      data_317 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_317 <= data_316;
        end
      end
    end
    if (reset) begin
      data_318 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_318 <= data_317;
        end
      end
    end
    if (reset) begin
      data_319 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_319 <= data_318;
        end
      end
    end
    if (reset) begin
      data_320 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_320 <= data_319;
        end
      end
    end
    if (reset) begin
      data_321 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_321 <= data_320;
        end
      end
    end
    if (reset) begin
      data_322 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_322 <= data_321;
        end
      end
    end
    if (reset) begin
      data_323 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_323 <= data_322;
        end
      end
    end
    if (reset) begin
      data_324 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_324 <= data_323;
        end
      end
    end
    if (reset) begin
      data_325 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_325 <= data_324;
        end
      end
    end
    if (reset) begin
      data_326 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_326 <= data_325;
        end
      end
    end
    if (reset) begin
      data_327 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_327 <= data_326;
        end
      end
    end
    if (reset) begin
      data_328 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_328 <= data_327;
        end
      end
    end
    if (reset) begin
      data_329 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_329 <= data_328;
        end
      end
    end
    if (reset) begin
      data_330 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_330 <= data_329;
        end
      end
    end
    if (reset) begin
      data_331 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_331 <= data_330;
        end
      end
    end
    if (reset) begin
      data_332 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_332 <= data_331;
        end
      end
    end
    if (reset) begin
      data_333 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_333 <= data_332;
        end
      end
    end
    if (reset) begin
      data_334 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_334 <= data_333;
        end
      end
    end
    if (reset) begin
      data_335 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_335 <= data_334;
        end
      end
    end
    if (reset) begin
      data_336 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_336 <= data_335;
        end
      end
    end
    if (reset) begin
      data_337 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_337 <= data_336;
        end
      end
    end
    if (reset) begin
      data_338 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_338 <= data_337;
        end
      end
    end
    if (reset) begin
      data_339 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_339 <= data_338;
        end
      end
    end
    if (reset) begin
      data_340 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_340 <= data_339;
        end
      end
    end
    if (reset) begin
      data_341 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_341 <= data_340;
        end
      end
    end
    if (reset) begin
      data_342 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_342 <= data_341;
        end
      end
    end
    if (reset) begin
      data_343 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_343 <= data_342;
        end
      end
    end
    if (reset) begin
      data_344 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_344 <= data_343;
        end
      end
    end
    if (reset) begin
      data_345 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_345 <= data_344;
        end
      end
    end
    if (reset) begin
      data_346 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_346 <= data_345;
        end
      end
    end
    if (reset) begin
      data_347 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_347 <= data_346;
        end
      end
    end
    if (reset) begin
      data_348 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_348 <= data_347;
        end
      end
    end
    if (reset) begin
      data_349 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_349 <= data_348;
        end
      end
    end
    if (reset) begin
      data_350 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_350 <= data_349;
        end
      end
    end
    if (reset) begin
      data_351 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_351 <= data_350;
        end
      end
    end
    if (reset) begin
      data_352 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_352 <= data_351;
        end
      end
    end
    if (reset) begin
      data_353 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_353 <= data_352;
        end
      end
    end
    if (reset) begin
      data_354 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_354 <= data_353;
        end
      end
    end
    if (reset) begin
      data_355 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_355 <= data_354;
        end
      end
    end
    if (reset) begin
      data_356 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_356 <= data_355;
        end
      end
    end
    if (reset) begin
      data_357 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_357 <= data_356;
        end
      end
    end
    if (reset) begin
      data_358 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_358 <= data_357;
        end
      end
    end
    if (reset) begin
      data_359 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_359 <= data_358;
        end
      end
    end
    if (reset) begin
      data_360 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_360 <= data_359;
        end
      end
    end
    if (reset) begin
      data_361 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_361 <= data_360;
        end
      end
    end
    if (reset) begin
      data_362 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_362 <= data_361;
        end
      end
    end
    if (reset) begin
      data_363 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_363 <= data_362;
        end
      end
    end
    if (reset) begin
      data_364 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_364 <= data_363;
        end
      end
    end
    if (reset) begin
      data_365 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_365 <= data_364;
        end
      end
    end
    if (reset) begin
      data_366 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_366 <= data_365;
        end
      end
    end
    if (reset) begin
      data_367 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_367 <= data_366;
        end
      end
    end
    if (reset) begin
      data_368 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_368 <= data_367;
        end
      end
    end
    if (reset) begin
      data_369 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_369 <= data_368;
        end
      end
    end
    if (reset) begin
      data_370 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_370 <= data_369;
        end
      end
    end
    if (reset) begin
      data_371 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_371 <= data_370;
        end
      end
    end
    if (reset) begin
      data_372 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_372 <= data_371;
        end
      end
    end
    if (reset) begin
      data_373 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_373 <= data_372;
        end
      end
    end
    if (reset) begin
      data_374 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_374 <= data_373;
        end
      end
    end
    if (reset) begin
      data_375 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_375 <= data_374;
        end
      end
    end
    if (reset) begin
      data_376 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_376 <= data_375;
        end
      end
    end
    if (reset) begin
      data_377 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_377 <= data_376;
        end
      end
    end
    if (reset) begin
      data_378 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_378 <= data_377;
        end
      end
    end
    if (reset) begin
      data_379 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_379 <= data_378;
        end
      end
    end
    if (reset) begin
      data_380 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_380 <= data_379;
        end
      end
    end
    if (reset) begin
      data_381 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_381 <= data_380;
        end
      end
    end
    if (reset) begin
      data_382 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_382 <= data_381;
        end
      end
    end
    if (reset) begin
      data_383 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_383 <= data_382;
        end
      end
    end
    if (reset) begin
      data_384 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_384 <= data_383;
        end
      end
    end
    if (reset) begin
      data_385 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_385 <= data_384;
        end
      end
    end
    if (reset) begin
      data_386 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_386 <= data_385;
        end
      end
    end
    if (reset) begin
      data_387 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_387 <= data_386;
        end
      end
    end
    if (reset) begin
      data_388 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_388 <= data_387;
        end
      end
    end
    if (reset) begin
      data_389 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_389 <= data_388;
        end
      end
    end
    if (reset) begin
      data_390 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_390 <= data_389;
        end
      end
    end
    if (reset) begin
      data_391 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_391 <= data_390;
        end
      end
    end
    if (reset) begin
      data_392 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_392 <= data_391;
        end
      end
    end
    if (reset) begin
      data_393 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_393 <= data_392;
        end
      end
    end
    if (reset) begin
      data_394 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_394 <= data_393;
        end
      end
    end
    if (reset) begin
      data_395 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_395 <= data_394;
        end
      end
    end
    if (reset) begin
      data_396 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_396 <= data_395;
        end
      end
    end
    if (reset) begin
      data_397 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_397 <= data_396;
        end
      end
    end
    if (reset) begin
      data_398 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_398 <= data_397;
        end
      end
    end
    if (reset) begin
      data_399 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_399 <= data_398;
        end
      end
    end
    if (reset) begin
      data_400 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_400 <= data_399;
        end
      end
    end
    if (reset) begin
      data_401 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_401 <= data_400;
        end
      end
    end
    if (reset) begin
      data_402 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_402 <= data_401;
        end
      end
    end
    if (reset) begin
      data_403 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_403 <= data_402;
        end
      end
    end
    if (reset) begin
      data_404 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_404 <= data_403;
        end
      end
    end
    if (reset) begin
      data_405 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_405 <= data_404;
        end
      end
    end
    if (reset) begin
      data_406 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_406 <= data_405;
        end
      end
    end
    if (reset) begin
      data_407 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_407 <= data_406;
        end
      end
    end
    if (reset) begin
      data_408 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_408 <= data_407;
        end
      end
    end
    if (reset) begin
      data_409 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_409 <= data_408;
        end
      end
    end
    if (reset) begin
      data_410 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_410 <= data_409;
        end
      end
    end
    if (reset) begin
      data_411 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_411 <= data_410;
        end
      end
    end
    if (reset) begin
      data_412 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_412 <= data_411;
        end
      end
    end
    if (reset) begin
      data_413 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_413 <= data_412;
        end
      end
    end
    if (reset) begin
      data_414 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_414 <= data_413;
        end
      end
    end
    if (reset) begin
      data_415 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_415 <= data_414;
        end
      end
    end
    if (reset) begin
      data_416 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_416 <= data_415;
        end
      end
    end
    if (reset) begin
      data_417 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_417 <= data_416;
        end
      end
    end
    if (reset) begin
      data_418 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_418 <= data_417;
        end
      end
    end
    if (reset) begin
      data_419 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_419 <= data_418;
        end
      end
    end
    if (reset) begin
      data_420 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_420 <= data_419;
        end
      end
    end
    if (reset) begin
      data_421 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_421 <= data_420;
        end
      end
    end
    if (reset) begin
      data_422 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_422 <= data_421;
        end
      end
    end
    if (reset) begin
      data_423 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_423 <= data_422;
        end
      end
    end
    if (reset) begin
      data_424 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_424 <= data_423;
        end
      end
    end
    if (reset) begin
      data_425 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_425 <= data_424;
        end
      end
    end
    if (reset) begin
      data_426 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_426 <= data_425;
        end
      end
    end
    if (reset) begin
      data_427 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_427 <= data_426;
        end
      end
    end
    if (reset) begin
      data_428 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_428 <= data_427;
        end
      end
    end
    if (reset) begin
      data_429 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_429 <= data_428;
        end
      end
    end
    if (reset) begin
      data_430 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_430 <= data_429;
        end
      end
    end
    if (reset) begin
      data_431 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_431 <= data_430;
        end
      end
    end
    if (reset) begin
      data_432 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_432 <= data_431;
        end
      end
    end
    if (reset) begin
      data_433 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_433 <= data_432;
        end
      end
    end
    if (reset) begin
      data_434 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_434 <= data_433;
        end
      end
    end
    if (reset) begin
      data_435 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_435 <= data_434;
        end
      end
    end
    if (reset) begin
      data_436 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_436 <= data_435;
        end
      end
    end
    if (reset) begin
      data_437 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_437 <= data_436;
        end
      end
    end
    if (reset) begin
      data_438 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_438 <= data_437;
        end
      end
    end
    if (reset) begin
      data_439 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_439 <= data_438;
        end
      end
    end
    if (reset) begin
      data_440 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_440 <= data_439;
        end
      end
    end
    if (reset) begin
      data_441 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_441 <= data_440;
        end
      end
    end
    if (reset) begin
      data_442 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_442 <= data_441;
        end
      end
    end
    if (reset) begin
      data_443 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_443 <= data_442;
        end
      end
    end
    if (reset) begin
      data_444 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_444 <= data_443;
        end
      end
    end
    if (reset) begin
      data_445 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_445 <= data_444;
        end
      end
    end
    if (reset) begin
      data_446 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_446 <= data_445;
        end
      end
    end
    if (reset) begin
      data_447 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_447 <= data_446;
        end
      end
    end
    if (reset) begin
      data_448 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_448 <= data_447;
        end
      end
    end
    if (reset) begin
      data_449 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_449 <= data_448;
        end
      end
    end
    if (reset) begin
      data_450 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_450 <= data_449;
        end
      end
    end
    if (reset) begin
      data_451 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_451 <= data_450;
        end
      end
    end
    if (reset) begin
      data_452 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_452 <= data_451;
        end
      end
    end
    if (reset) begin
      data_453 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_453 <= data_452;
        end
      end
    end
    if (reset) begin
      data_454 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_454 <= data_453;
        end
      end
    end
    if (reset) begin
      data_455 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_455 <= data_454;
        end
      end
    end
    if (reset) begin
      data_456 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_456 <= data_455;
        end
      end
    end
    if (reset) begin
      data_457 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_457 <= data_456;
        end
      end
    end
    if (reset) begin
      data_458 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_458 <= data_457;
        end
      end
    end
    if (reset) begin
      data_459 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_459 <= data_458;
        end
      end
    end
    if (reset) begin
      data_460 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_460 <= data_459;
        end
      end
    end
    if (reset) begin
      data_461 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_461 <= data_460;
        end
      end
    end
    if (reset) begin
      data_462 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_462 <= data_461;
        end
      end
    end
    if (reset) begin
      data_463 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_463 <= data_462;
        end
      end
    end
    if (reset) begin
      data_464 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_464 <= data_463;
        end
      end
    end
    if (reset) begin
      data_465 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_465 <= data_464;
        end
      end
    end
    if (reset) begin
      data_466 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_466 <= data_465;
        end
      end
    end
    if (reset) begin
      data_467 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_467 <= data_466;
        end
      end
    end
    if (reset) begin
      data_468 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_468 <= data_467;
        end
      end
    end
    if (reset) begin
      data_469 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_469 <= data_468;
        end
      end
    end
    if (reset) begin
      data_470 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_470 <= data_469;
        end
      end
    end
    if (reset) begin
      data_471 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_471 <= data_470;
        end
      end
    end
    if (reset) begin
      data_472 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_472 <= data_471;
        end
      end
    end
    if (reset) begin
      data_473 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_473 <= data_472;
        end
      end
    end
    if (reset) begin
      data_474 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_474 <= data_473;
        end
      end
    end
    if (reset) begin
      data_475 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_475 <= data_474;
        end
      end
    end
    if (reset) begin
      data_476 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_476 <= data_475;
        end
      end
    end
    if (reset) begin
      data_477 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_477 <= data_476;
        end
      end
    end
    if (reset) begin
      data_478 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_478 <= data_477;
        end
      end
    end
    if (reset) begin
      data_479 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_479 <= data_478;
        end
      end
    end
    if (reset) begin
      data_480 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_480 <= data_479;
        end
      end
    end
    if (reset) begin
      data_481 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_481 <= data_480;
        end
      end
    end
    if (reset) begin
      data_482 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_482 <= data_481;
        end
      end
    end
    if (reset) begin
      data_483 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_483 <= data_482;
        end
      end
    end
    if (reset) begin
      data_484 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_484 <= data_483;
        end
      end
    end
    if (reset) begin
      data_485 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_485 <= data_484;
        end
      end
    end
    if (reset) begin
      data_486 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_486 <= data_485;
        end
      end
    end
    if (reset) begin
      data_487 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_487 <= data_486;
        end
      end
    end
    if (reset) begin
      data_488 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_488 <= data_487;
        end
      end
    end
    if (reset) begin
      data_489 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_489 <= data_488;
        end
      end
    end
    if (reset) begin
      data_490 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_490 <= data_489;
        end
      end
    end
    if (reset) begin
      data_491 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_491 <= data_490;
        end
      end
    end
    if (reset) begin
      data_492 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_492 <= data_491;
        end
      end
    end
    if (reset) begin
      data_493 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_493 <= data_492;
        end
      end
    end
    if (reset) begin
      data_494 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_494 <= data_493;
        end
      end
    end
    if (reset) begin
      data_495 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_495 <= data_494;
        end
      end
    end
    if (reset) begin
      data_496 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_496 <= data_495;
        end
      end
    end
    if (reset) begin
      data_497 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_497 <= data_496;
        end
      end
    end
    if (reset) begin
      data_498 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_498 <= data_497;
        end
      end
    end
    if (reset) begin
      data_499 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_499 <= data_498;
        end
      end
    end
    if (reset) begin
      data_500 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_500 <= data_499;
        end
      end
    end
    if (reset) begin
      data_501 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_501 <= data_500;
        end
      end
    end
    if (reset) begin
      data_502 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_502 <= data_501;
        end
      end
    end
    if (reset) begin
      data_503 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_503 <= data_502;
        end
      end
    end
    if (reset) begin
      data_504 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_504 <= data_503;
        end
      end
    end
    if (reset) begin
      data_505 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_505 <= data_504;
        end
      end
    end
    if (reset) begin
      data_506 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_506 <= data_505;
        end
      end
    end
    if (reset) begin
      data_507 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_507 <= data_506;
        end
      end
    end
    if (reset) begin
      data_508 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_508 <= data_507;
        end
      end
    end
    if (reset) begin
      data_509 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_509 <= data_508;
        end
      end
    end
    if (reset) begin
      data_510 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_510 <= data_509;
        end
      end
    end
    if (reset) begin
      data_511 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_511 <= data_510;
        end
      end
    end
    if (reset) begin
      data_512 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_512 <= data_511;
        end
      end
    end
    if (reset) begin
      data_513 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_513 <= data_512;
        end
      end
    end
    if (reset) begin
      data_514 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_514 <= data_513;
        end
      end
    end
    if (reset) begin
      data_515 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_515 <= data_514;
        end
      end
    end
    if (reset) begin
      data_516 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_516 <= data_515;
        end
      end
    end
    if (reset) begin
      data_517 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_517 <= data_516;
        end
      end
    end
    if (reset) begin
      data_518 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_518 <= data_517;
        end
      end
    end
    if (reset) begin
      data_519 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_519 <= data_518;
        end
      end
    end
    if (reset) begin
      data_520 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_520 <= data_519;
        end
      end
    end
    if (reset) begin
      data_521 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_521 <= data_520;
        end
      end
    end
    if (reset) begin
      data_522 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_522 <= data_521;
        end
      end
    end
    if (reset) begin
      data_523 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_523 <= data_522;
        end
      end
    end
    if (reset) begin
      data_524 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_524 <= data_523;
        end
      end
    end
    if (reset) begin
      data_525 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_525 <= data_524;
        end
      end
    end
    if (reset) begin
      data_526 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_526 <= data_525;
        end
      end
    end
    if (reset) begin
      data_527 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_527 <= data_526;
        end
      end
    end
    if (reset) begin
      data_528 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_528 <= data_527;
        end
      end
    end
    if (reset) begin
      data_529 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_529 <= data_528;
        end
      end
    end
    if (reset) begin
      data_530 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_530 <= data_529;
        end
      end
    end
    if (reset) begin
      data_531 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_531 <= data_530;
        end
      end
    end
    if (reset) begin
      data_532 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_532 <= data_531;
        end
      end
    end
    if (reset) begin
      data_533 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_533 <= data_532;
        end
      end
    end
    if (reset) begin
      data_534 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_534 <= data_533;
        end
      end
    end
    if (reset) begin
      data_535 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_535 <= data_534;
        end
      end
    end
    if (reset) begin
      data_536 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_536 <= data_535;
        end
      end
    end
    if (reset) begin
      data_537 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_537 <= data_536;
        end
      end
    end
    if (reset) begin
      data_538 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_538 <= data_537;
        end
      end
    end
    if (reset) begin
      data_539 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_539 <= data_538;
        end
      end
    end
    if (reset) begin
      data_540 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_540 <= data_539;
        end
      end
    end
    if (reset) begin
      data_541 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_541 <= data_540;
        end
      end
    end
    if (reset) begin
      data_542 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_542 <= data_541;
        end
      end
    end
    if (reset) begin
      data_543 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_543 <= data_542;
        end
      end
    end
    if (reset) begin
      data_544 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_544 <= data_543;
        end
      end
    end
    if (reset) begin
      data_545 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_545 <= data_544;
        end
      end
    end
    if (reset) begin
      data_546 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_546 <= data_545;
        end
      end
    end
    if (reset) begin
      data_547 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_547 <= data_546;
        end
      end
    end
    if (reset) begin
      data_548 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_548 <= data_547;
        end
      end
    end
    if (reset) begin
      data_549 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_549 <= data_548;
        end
      end
    end
    if (reset) begin
      data_550 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_550 <= data_549;
        end
      end
    end
    if (reset) begin
      data_551 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_551 <= data_550;
        end
      end
    end
    if (reset) begin
      data_552 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_552 <= data_551;
        end
      end
    end
    if (reset) begin
      data_553 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_553 <= data_552;
        end
      end
    end
    if (reset) begin
      data_554 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_554 <= data_553;
        end
      end
    end
    if (reset) begin
      data_555 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_555 <= data_554;
        end
      end
    end
    if (reset) begin
      data_556 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_556 <= data_555;
        end
      end
    end
    if (reset) begin
      data_557 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_557 <= data_556;
        end
      end
    end
    if (reset) begin
      data_558 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_558 <= data_557;
        end
      end
    end
    if (reset) begin
      data_559 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_559 <= data_558;
        end
      end
    end
    if (reset) begin
      data_560 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_560 <= data_559;
        end
      end
    end
    if (reset) begin
      data_561 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_561 <= data_560;
        end
      end
    end
    if (reset) begin
      data_562 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_562 <= data_561;
        end
      end
    end
    if (reset) begin
      data_563 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_563 <= data_562;
        end
      end
    end
    if (reset) begin
      data_564 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_564 <= data_563;
        end
      end
    end
    if (reset) begin
      data_565 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_565 <= data_564;
        end
      end
    end
    if (reset) begin
      data_566 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_566 <= data_565;
        end
      end
    end
    if (reset) begin
      data_567 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_567 <= data_566;
        end
      end
    end
    if (reset) begin
      data_568 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_568 <= data_567;
        end
      end
    end
    if (reset) begin
      data_569 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_569 <= data_568;
        end
      end
    end
    if (reset) begin
      data_570 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_570 <= data_569;
        end
      end
    end
    if (reset) begin
      data_571 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_571 <= data_570;
        end
      end
    end
    if (reset) begin
      data_572 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_572 <= data_571;
        end
      end
    end
    if (reset) begin
      data_573 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_573 <= data_572;
        end
      end
    end
    if (reset) begin
      data_574 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_574 <= data_573;
        end
      end
    end
    if (reset) begin
      data_575 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_575 <= data_574;
        end
      end
    end
    if (reset) begin
      data_576 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_576 <= data_575;
        end
      end
    end
    if (reset) begin
      data_577 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_577 <= data_576;
        end
      end
    end
    if (reset) begin
      data_578 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_578 <= data_577;
        end
      end
    end
    if (reset) begin
      data_579 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_579 <= data_578;
        end
      end
    end
    if (reset) begin
      data_580 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_580 <= data_579;
        end
      end
    end
    if (reset) begin
      data_581 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_581 <= data_580;
        end
      end
    end
    if (reset) begin
      data_582 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_582 <= data_581;
        end
      end
    end
    if (reset) begin
      data_583 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_583 <= data_582;
        end
      end
    end
    if (reset) begin
      data_584 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_584 <= data_583;
        end
      end
    end
    if (reset) begin
      data_585 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_585 <= data_584;
        end
      end
    end
    if (reset) begin
      data_586 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_586 <= data_585;
        end
      end
    end
    if (reset) begin
      data_587 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_587 <= data_586;
        end
      end
    end
    if (reset) begin
      data_588 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_588 <= data_587;
        end
      end
    end
    if (reset) begin
      data_589 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_589 <= data_588;
        end
      end
    end
    if (reset) begin
      data_590 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_590 <= data_589;
        end
      end
    end
    if (reset) begin
      data_591 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_591 <= data_590;
        end
      end
    end
    if (reset) begin
      data_592 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_592 <= data_591;
        end
      end
    end
    if (reset) begin
      data_593 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_593 <= data_592;
        end
      end
    end
    if (reset) begin
      data_594 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_594 <= data_593;
        end
      end
    end
    if (reset) begin
      data_595 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_595 <= data_594;
        end
      end
    end
    if (reset) begin
      data_596 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_596 <= data_595;
        end
      end
    end
    if (reset) begin
      data_597 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_597 <= data_596;
        end
      end
    end
    if (reset) begin
      data_598 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_598 <= data_597;
        end
      end
    end
    if (reset) begin
      data_599 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_599 <= data_598;
        end
      end
    end
    if (reset) begin
      data_600 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_600 <= data_599;
        end
      end
    end
    if (reset) begin
      data_601 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_601 <= data_600;
        end
      end
    end
    if (reset) begin
      data_602 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_602 <= data_601;
        end
      end
    end
    if (reset) begin
      data_603 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_603 <= data_602;
        end
      end
    end
    if (reset) begin
      data_604 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_604 <= data_603;
        end
      end
    end
    if (reset) begin
      data_605 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_605 <= data_604;
        end
      end
    end
    if (reset) begin
      data_606 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_606 <= data_605;
        end
      end
    end
    if (reset) begin
      data_607 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_607 <= data_606;
        end
      end
    end
    if (reset) begin
      data_608 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_608 <= data_607;
        end
      end
    end
    if (reset) begin
      data_609 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_609 <= data_608;
        end
      end
    end
    if (reset) begin
      data_610 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_610 <= data_609;
        end
      end
    end
    if (reset) begin
      data_611 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_611 <= data_610;
        end
      end
    end
    if (reset) begin
      data_612 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_612 <= data_611;
        end
      end
    end
    if (reset) begin
      data_613 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_613 <= data_612;
        end
      end
    end
    if (reset) begin
      data_614 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_614 <= data_613;
        end
      end
    end
    if (reset) begin
      data_615 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_615 <= data_614;
        end
      end
    end
    if (reset) begin
      data_616 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_616 <= data_615;
        end
      end
    end
    if (reset) begin
      data_617 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_617 <= data_616;
        end
      end
    end
    if (reset) begin
      data_618 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_618 <= data_617;
        end
      end
    end
    if (reset) begin
      data_619 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_619 <= data_618;
        end
      end
    end
    if (reset) begin
      data_620 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_620 <= data_619;
        end
      end
    end
    if (reset) begin
      data_621 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_621 <= data_620;
        end
      end
    end
    if (reset) begin
      data_622 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_622 <= data_621;
        end
      end
    end
    if (reset) begin
      data_623 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_623 <= data_622;
        end
      end
    end
    if (reset) begin
      data_624 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_624 <= data_623;
        end
      end
    end
    if (reset) begin
      data_625 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_625 <= data_624;
        end
      end
    end
    if (reset) begin
      data_626 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_626 <= data_625;
        end
      end
    end
    if (reset) begin
      data_627 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_627 <= data_626;
        end
      end
    end
    if (reset) begin
      data_628 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_628 <= data_627;
        end
      end
    end
    if (reset) begin
      data_629 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_629 <= data_628;
        end
      end
    end
    if (reset) begin
      data_630 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_630 <= data_629;
        end
      end
    end
    if (reset) begin
      data_631 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_631 <= data_630;
        end
      end
    end
    if (reset) begin
      data_632 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_632 <= data_631;
        end
      end
    end
    if (reset) begin
      data_633 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_633 <= data_632;
        end
      end
    end
    if (reset) begin
      data_634 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_634 <= data_633;
        end
      end
    end
    if (reset) begin
      data_635 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_635 <= data_634;
        end
      end
    end
    if (reset) begin
      data_636 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_636 <= data_635;
        end
      end
    end
    if (reset) begin
      data_637 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_637 <= data_636;
        end
      end
    end
    if (reset) begin
      data_638 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_638 <= data_637;
        end
      end
    end
    if (reset) begin
      data_639 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_639 <= data_638;
        end
      end
    end
    if (reset) begin
      data_640 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_640 <= data_639;
        end
      end
    end
    if (reset) begin
      data_641 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_641 <= data_640;
        end
      end
    end
    if (reset) begin
      data_642 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_642 <= data_641;
        end
      end
    end
    if (reset) begin
      data_643 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_643 <= data_642;
        end
      end
    end
    if (reset) begin
      data_644 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_644 <= data_643;
        end
      end
    end
    if (reset) begin
      data_645 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_645 <= data_644;
        end
      end
    end
    if (reset) begin
      data_646 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_646 <= data_645;
        end
      end
    end
    if (reset) begin
      data_647 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_647 <= data_646;
        end
      end
    end
    if (reset) begin
      data_648 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_648 <= data_647;
        end
      end
    end
    if (reset) begin
      data_649 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_649 <= data_648;
        end
      end
    end
    if (reset) begin
      data_650 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_650 <= data_649;
        end
      end
    end
    if (reset) begin
      data_651 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_651 <= data_650;
        end
      end
    end
    if (reset) begin
      data_652 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_652 <= data_651;
        end
      end
    end
    if (reset) begin
      data_653 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_653 <= data_652;
        end
      end
    end
    if (reset) begin
      data_654 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_654 <= data_653;
        end
      end
    end
    if (reset) begin
      data_655 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_655 <= data_654;
        end
      end
    end
    if (reset) begin
      data_656 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_656 <= data_655;
        end
      end
    end
    if (reset) begin
      data_657 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_657 <= data_656;
        end
      end
    end
    if (reset) begin
      data_658 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_658 <= data_657;
        end
      end
    end
    if (reset) begin
      data_659 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_659 <= data_658;
        end
      end
    end
    if (reset) begin
      data_660 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_660 <= data_659;
        end
      end
    end
    if (reset) begin
      data_661 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_661 <= data_660;
        end
      end
    end
    if (reset) begin
      data_662 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_662 <= data_661;
        end
      end
    end
    if (reset) begin
      data_663 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_663 <= data_662;
        end
      end
    end
    if (reset) begin
      data_664 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_664 <= data_663;
        end
      end
    end
    if (reset) begin
      data_665 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_665 <= data_664;
        end
      end
    end
    if (reset) begin
      data_666 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_666 <= data_665;
        end
      end
    end
    if (reset) begin
      data_667 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_667 <= data_666;
        end
      end
    end
    if (reset) begin
      data_668 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_668 <= data_667;
        end
      end
    end
    if (reset) begin
      data_669 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_669 <= data_668;
        end
      end
    end
    if (reset) begin
      data_670 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_670 <= data_669;
        end
      end
    end
    if (reset) begin
      data_671 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_671 <= data_670;
        end
      end
    end
    if (reset) begin
      data_672 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_672 <= data_671;
        end
      end
    end
    if (reset) begin
      data_673 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_673 <= data_672;
        end
      end
    end
    if (reset) begin
      data_674 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_674 <= data_673;
        end
      end
    end
    if (reset) begin
      data_675 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_675 <= data_674;
        end
      end
    end
    if (reset) begin
      data_676 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_676 <= data_675;
        end
      end
    end
    if (reset) begin
      data_677 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_677 <= data_676;
        end
      end
    end
    if (reset) begin
      data_678 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_678 <= data_677;
        end
      end
    end
    if (reset) begin
      data_679 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_679 <= data_678;
        end
      end
    end
    if (reset) begin
      data_680 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_680 <= data_679;
        end
      end
    end
    if (reset) begin
      data_681 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_681 <= data_680;
        end
      end
    end
    if (reset) begin
      data_682 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_682 <= data_681;
        end
      end
    end
    if (reset) begin
      data_683 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_683 <= data_682;
        end
      end
    end
    if (reset) begin
      data_684 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_684 <= data_683;
        end
      end
    end
    if (reset) begin
      data_685 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_685 <= data_684;
        end
      end
    end
    if (reset) begin
      data_686 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_686 <= data_685;
        end
      end
    end
    if (reset) begin
      data_687 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_687 <= data_686;
        end
      end
    end
    if (reset) begin
      data_688 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_688 <= data_687;
        end
      end
    end
    if (reset) begin
      data_689 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_689 <= data_688;
        end
      end
    end
    if (reset) begin
      data_690 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_690 <= data_689;
        end
      end
    end
    if (reset) begin
      data_691 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_691 <= data_690;
        end
      end
    end
    if (reset) begin
      data_692 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_692 <= data_691;
        end
      end
    end
    if (reset) begin
      data_693 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_693 <= data_692;
        end
      end
    end
    if (reset) begin
      data_694 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_694 <= data_693;
        end
      end
    end
    if (reset) begin
      data_695 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_695 <= data_694;
        end
      end
    end
    if (reset) begin
      data_696 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_696 <= data_695;
        end
      end
    end
    if (reset) begin
      data_697 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_697 <= data_696;
        end
      end
    end
    if (reset) begin
      data_698 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_698 <= data_697;
        end
      end
    end
    if (reset) begin
      data_699 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_699 <= data_698;
        end
      end
    end
    if (reset) begin
      data_700 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_700 <= data_699;
        end
      end
    end
    if (reset) begin
      data_701 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_701 <= data_700;
        end
      end
    end
    if (reset) begin
      data_702 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_702 <= data_701;
        end
      end
    end
    if (reset) begin
      data_703 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_703 <= data_702;
        end
      end
    end
    if (reset) begin
      data_704 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_704 <= data_703;
        end
      end
    end
    if (reset) begin
      data_705 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_705 <= data_704;
        end
      end
    end
    if (reset) begin
      data_706 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_706 <= data_705;
        end
      end
    end
    if (reset) begin
      data_707 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_707 <= data_706;
        end
      end
    end
    if (reset) begin
      data_708 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_708 <= data_707;
        end
      end
    end
    if (reset) begin
      data_709 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_709 <= data_708;
        end
      end
    end
    if (reset) begin
      data_710 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_710 <= data_709;
        end
      end
    end
    if (reset) begin
      data_711 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_711 <= data_710;
        end
      end
    end
    if (reset) begin
      data_712 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_712 <= data_711;
        end
      end
    end
    if (reset) begin
      data_713 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_713 <= data_712;
        end
      end
    end
    if (reset) begin
      data_714 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_714 <= data_713;
        end
      end
    end
    if (reset) begin
      data_715 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_715 <= data_714;
        end
      end
    end
    if (reset) begin
      data_716 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_716 <= data_715;
        end
      end
    end
    if (reset) begin
      data_717 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_717 <= data_716;
        end
      end
    end
    if (reset) begin
      data_718 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_718 <= data_717;
        end
      end
    end
    if (reset) begin
      data_719 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_719 <= data_718;
        end
      end
    end
    if (reset) begin
      data_720 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_720 <= data_719;
        end
      end
    end
    if (reset) begin
      data_721 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_721 <= data_720;
        end
      end
    end
    if (reset) begin
      data_722 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_722 <= data_721;
        end
      end
    end
    if (reset) begin
      data_723 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_723 <= data_722;
        end
      end
    end
    if (reset) begin
      data_724 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_724 <= data_723;
        end
      end
    end
    if (reset) begin
      data_725 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_725 <= data_724;
        end
      end
    end
    if (reset) begin
      data_726 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_726 <= data_725;
        end
      end
    end
    if (reset) begin
      data_727 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_727 <= data_726;
        end
      end
    end
    if (reset) begin
      data_728 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_728 <= data_727;
        end
      end
    end
    if (reset) begin
      data_729 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_729 <= data_728;
        end
      end
    end
    if (reset) begin
      data_730 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_730 <= data_729;
        end
      end
    end
    if (reset) begin
      data_731 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_731 <= data_730;
        end
      end
    end
    if (reset) begin
      data_732 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_732 <= data_731;
        end
      end
    end
    if (reset) begin
      data_733 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_733 <= data_732;
        end
      end
    end
    if (reset) begin
      data_734 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_734 <= data_733;
        end
      end
    end
    if (reset) begin
      data_735 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_735 <= data_734;
        end
      end
    end
    if (reset) begin
      data_736 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_736 <= data_735;
        end
      end
    end
    if (reset) begin
      data_737 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_737 <= data_736;
        end
      end
    end
    if (reset) begin
      data_738 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_738 <= data_737;
        end
      end
    end
    if (reset) begin
      data_739 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_739 <= data_738;
        end
      end
    end
    if (reset) begin
      data_740 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_740 <= data_739;
        end
      end
    end
    if (reset) begin
      data_741 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_741 <= data_740;
        end
      end
    end
    if (reset) begin
      data_742 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_742 <= data_741;
        end
      end
    end
    if (reset) begin
      data_743 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_743 <= data_742;
        end
      end
    end
    if (reset) begin
      data_744 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_744 <= data_743;
        end
      end
    end
    if (reset) begin
      data_745 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_745 <= data_744;
        end
      end
    end
    if (reset) begin
      data_746 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_746 <= data_745;
        end
      end
    end
    if (reset) begin
      data_747 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_747 <= data_746;
        end
      end
    end
    if (reset) begin
      data_748 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_748 <= data_747;
        end
      end
    end
    if (reset) begin
      data_749 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_749 <= data_748;
        end
      end
    end
    if (reset) begin
      data_750 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_750 <= data_749;
        end
      end
    end
    if (reset) begin
      data_751 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_751 <= data_750;
        end
      end
    end
    if (reset) begin
      data_752 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_752 <= data_751;
        end
      end
    end
    if (reset) begin
      data_753 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_753 <= data_752;
        end
      end
    end
    if (reset) begin
      data_754 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_754 <= data_753;
        end
      end
    end
    if (reset) begin
      data_755 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_755 <= data_754;
        end
      end
    end
    if (reset) begin
      data_756 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_756 <= data_755;
        end
      end
    end
    if (reset) begin
      data_757 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_757 <= data_756;
        end
      end
    end
    if (reset) begin
      data_758 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_758 <= data_757;
        end
      end
    end
    if (reset) begin
      data_759 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_759 <= data_758;
        end
      end
    end
    if (reset) begin
      data_760 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_760 <= data_759;
        end
      end
    end
    if (reset) begin
      data_761 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_761 <= data_760;
        end
      end
    end
    if (reset) begin
      data_762 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_762 <= data_761;
        end
      end
    end
    if (reset) begin
      data_763 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_763 <= data_762;
        end
      end
    end
    if (reset) begin
      data_764 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_764 <= data_763;
        end
      end
    end
    if (reset) begin
      data_765 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_765 <= data_764;
        end
      end
    end
    if (reset) begin
      data_766 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_766 <= data_765;
        end
      end
    end
    if (reset) begin
      data_767 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_767 <= data_766;
        end
      end
    end
    if (reset) begin
      data_768 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_768 <= data_767;
        end
      end
    end
    if (reset) begin
      data_769 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_769 <= data_768;
        end
      end
    end
    if (reset) begin
      data_770 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_770 <= data_769;
        end
      end
    end
    if (reset) begin
      data_771 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_771 <= data_770;
        end
      end
    end
    if (reset) begin
      data_772 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_772 <= data_771;
        end
      end
    end
    if (reset) begin
      data_773 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_773 <= data_772;
        end
      end
    end
    if (reset) begin
      data_774 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_774 <= data_773;
        end
      end
    end
    if (reset) begin
      data_775 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_775 <= data_774;
        end
      end
    end
    if (reset) begin
      data_776 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_776 <= data_775;
        end
      end
    end
    if (reset) begin
      data_777 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_777 <= data_776;
        end
      end
    end
    if (reset) begin
      data_778 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_778 <= data_777;
        end
      end
    end
    if (reset) begin
      data_779 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_779 <= data_778;
        end
      end
    end
    if (reset) begin
      data_780 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_780 <= data_779;
        end
      end
    end
    if (reset) begin
      data_781 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_781 <= data_780;
        end
      end
    end
    if (reset) begin
      data_782 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_782 <= data_781;
        end
      end
    end
    if (reset) begin
      data_783 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_783 <= data_782;
        end
      end
    end
    if (reset) begin
      data_784 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_784 <= data_783;
        end
      end
    end
    if (reset) begin
      data_785 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_785 <= data_784;
        end
      end
    end
    if (reset) begin
      data_786 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_786 <= data_785;
        end
      end
    end
    if (reset) begin
      data_787 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_787 <= data_786;
        end
      end
    end
    if (reset) begin
      data_788 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_788 <= data_787;
        end
      end
    end
    if (reset) begin
      data_789 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_789 <= data_788;
        end
      end
    end
    if (reset) begin
      data_790 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_790 <= data_789;
        end
      end
    end
    if (reset) begin
      data_791 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_791 <= data_790;
        end
      end
    end
    if (reset) begin
      data_792 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_792 <= data_791;
        end
      end
    end
    if (reset) begin
      data_793 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_793 <= data_792;
        end
      end
    end
    if (reset) begin
      data_794 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_794 <= data_793;
        end
      end
    end
    if (reset) begin
      data_795 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_795 <= data_794;
        end
      end
    end
    if (reset) begin
      data_796 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_796 <= data_795;
        end
      end
    end
    if (reset) begin
      data_797 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_797 <= data_796;
        end
      end
    end
    if (reset) begin
      data_798 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_798 <= data_797;
        end
      end
    end
    if (reset) begin
      data_799 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_799 <= data_798;
        end
      end
    end
    if (reset) begin
      data_800 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_800 <= data_799;
        end
      end
    end
    if (reset) begin
      data_801 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_801 <= data_800;
        end
      end
    end
    if (reset) begin
      data_802 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_802 <= data_801;
        end
      end
    end
    if (reset) begin
      data_803 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_803 <= data_802;
        end
      end
    end
    if (reset) begin
      data_804 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_804 <= data_803;
        end
      end
    end
    if (reset) begin
      data_805 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_805 <= data_804;
        end
      end
    end
    if (reset) begin
      data_806 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_806 <= data_805;
        end
      end
    end
    if (reset) begin
      data_807 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_807 <= data_806;
        end
      end
    end
    if (reset) begin
      data_808 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_808 <= data_807;
        end
      end
    end
    if (reset) begin
      data_809 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_809 <= data_808;
        end
      end
    end
    if (reset) begin
      data_810 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_810 <= data_809;
        end
      end
    end
    if (reset) begin
      data_811 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_811 <= data_810;
        end
      end
    end
    if (reset) begin
      data_812 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_812 <= data_811;
        end
      end
    end
    if (reset) begin
      data_813 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_813 <= data_812;
        end
      end
    end
    if (reset) begin
      data_814 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_814 <= data_813;
        end
      end
    end
    if (reset) begin
      data_815 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_815 <= data_814;
        end
      end
    end
    if (reset) begin
      data_816 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_816 <= data_815;
        end
      end
    end
    if (reset) begin
      data_817 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_817 <= data_816;
        end
      end
    end
    if (reset) begin
      data_818 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_818 <= data_817;
        end
      end
    end
    if (reset) begin
      data_819 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_819 <= data_818;
        end
      end
    end
    if (reset) begin
      data_820 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_820 <= data_819;
        end
      end
    end
    if (reset) begin
      data_821 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_821 <= data_820;
        end
      end
    end
    if (reset) begin
      data_822 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_822 <= data_821;
        end
      end
    end
    if (reset) begin
      data_823 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_823 <= data_822;
        end
      end
    end
    if (reset) begin
      data_824 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_824 <= data_823;
        end
      end
    end
    if (reset) begin
      data_825 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_825 <= data_824;
        end
      end
    end
    if (reset) begin
      data_826 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_826 <= data_825;
        end
      end
    end
    if (reset) begin
      data_827 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_827 <= data_826;
        end
      end
    end
    if (reset) begin
      data_828 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_828 <= data_827;
        end
      end
    end
    if (reset) begin
      data_829 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_829 <= data_828;
        end
      end
    end
    if (reset) begin
      data_830 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_830 <= data_829;
        end
      end
    end
    if (reset) begin
      data_831 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_831 <= data_830;
        end
      end
    end
    if (reset) begin
      data_832 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_832 <= data_831;
        end
      end
    end
    if (reset) begin
      data_833 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_833 <= data_832;
        end
      end
    end
    if (reset) begin
      data_834 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_834 <= data_833;
        end
      end
    end
    if (reset) begin
      data_835 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_835 <= data_834;
        end
      end
    end
    if (reset) begin
      data_836 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_836 <= data_835;
        end
      end
    end
    if (reset) begin
      data_837 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_837 <= data_836;
        end
      end
    end
    if (reset) begin
      data_838 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_838 <= data_837;
        end
      end
    end
    if (reset) begin
      data_839 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_839 <= data_838;
        end
      end
    end
    if (reset) begin
      data_840 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_840 <= data_839;
        end
      end
    end
    if (reset) begin
      data_841 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_841 <= data_840;
        end
      end
    end
    if (reset) begin
      data_842 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_842 <= data_841;
        end
      end
    end
    if (reset) begin
      data_843 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_843 <= data_842;
        end
      end
    end
    if (reset) begin
      data_844 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_844 <= data_843;
        end
      end
    end
    if (reset) begin
      data_845 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_845 <= data_844;
        end
      end
    end
    if (reset) begin
      data_846 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_846 <= data_845;
        end
      end
    end
    if (reset) begin
      data_847 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_847 <= data_846;
        end
      end
    end
    if (reset) begin
      data_848 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_848 <= data_847;
        end
      end
    end
    if (reset) begin
      data_849 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_849 <= data_848;
        end
      end
    end
    if (reset) begin
      data_850 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_850 <= data_849;
        end
      end
    end
    if (reset) begin
      data_851 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_851 <= data_850;
        end
      end
    end
    if (reset) begin
      data_852 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_852 <= data_851;
        end
      end
    end
    if (reset) begin
      data_853 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_853 <= data_852;
        end
      end
    end
    if (reset) begin
      data_854 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_854 <= data_853;
        end
      end
    end
    if (reset) begin
      data_855 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_855 <= data_854;
        end
      end
    end
    if (reset) begin
      data_856 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_856 <= data_855;
        end
      end
    end
    if (reset) begin
      data_857 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_857 <= data_856;
        end
      end
    end
    if (reset) begin
      data_858 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_858 <= data_857;
        end
      end
    end
    if (reset) begin
      data_859 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_859 <= data_858;
        end
      end
    end
    if (reset) begin
      data_860 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_860 <= data_859;
        end
      end
    end
    if (reset) begin
      data_861 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_861 <= data_860;
        end
      end
    end
    if (reset) begin
      data_862 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_862 <= data_861;
        end
      end
    end
    if (reset) begin
      data_863 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_863 <= data_862;
        end
      end
    end
    if (reset) begin
      data_864 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_864 <= data_863;
        end
      end
    end
    if (reset) begin
      data_865 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_865 <= data_864;
        end
      end
    end
    if (reset) begin
      data_866 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_866 <= data_865;
        end
      end
    end
    if (reset) begin
      data_867 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_867 <= data_866;
        end
      end
    end
    if (reset) begin
      data_868 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_868 <= data_867;
        end
      end
    end
    if (reset) begin
      data_869 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_869 <= data_868;
        end
      end
    end
    if (reset) begin
      data_870 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_870 <= data_869;
        end
      end
    end
    if (reset) begin
      data_871 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_871 <= data_870;
        end
      end
    end
    if (reset) begin
      data_872 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_872 <= data_871;
        end
      end
    end
    if (reset) begin
      data_873 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_873 <= data_872;
        end
      end
    end
    if (reset) begin
      data_874 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_874 <= data_873;
        end
      end
    end
    if (reset) begin
      data_875 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_875 <= data_874;
        end
      end
    end
    if (reset) begin
      data_876 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_876 <= data_875;
        end
      end
    end
    if (reset) begin
      data_877 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_877 <= data_876;
        end
      end
    end
    if (reset) begin
      data_878 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_878 <= data_877;
        end
      end
    end
    if (reset) begin
      data_879 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_879 <= data_878;
        end
      end
    end
    if (reset) begin
      data_880 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_880 <= data_879;
        end
      end
    end
    if (reset) begin
      data_881 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_881 <= data_880;
        end
      end
    end
    if (reset) begin
      data_882 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_882 <= data_881;
        end
      end
    end
    if (reset) begin
      data_883 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_883 <= data_882;
        end
      end
    end
    if (reset) begin
      data_884 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_884 <= data_883;
        end
      end
    end
    if (reset) begin
      data_885 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_885 <= data_884;
        end
      end
    end
    if (reset) begin
      data_886 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_886 <= data_885;
        end
      end
    end
    if (reset) begin
      data_887 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_887 <= data_886;
        end
      end
    end
    if (reset) begin
      data_888 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_888 <= data_887;
        end
      end
    end
    if (reset) begin
      data_889 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_889 <= data_888;
        end
      end
    end
    if (reset) begin
      data_890 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_890 <= data_889;
        end
      end
    end
    if (reset) begin
      data_891 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_891 <= data_890;
        end
      end
    end
    if (reset) begin
      data_892 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_892 <= data_891;
        end
      end
    end
    if (reset) begin
      data_893 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_893 <= data_892;
        end
      end
    end
    if (reset) begin
      data_894 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_894 <= data_893;
        end
      end
    end
    if (reset) begin
      data_895 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_895 <= data_894;
        end
      end
    end
    if (reset) begin
      data_896 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_896 <= data_895;
        end
      end
    end
    if (reset) begin
      data_897 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_897 <= data_896;
        end
      end
    end
    if (reset) begin
      data_898 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_898 <= data_897;
        end
      end
    end
    if (reset) begin
      data_899 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_899 <= data_898;
        end
      end
    end
    if (reset) begin
      data_900 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_900 <= data_899;
        end
      end
    end
    if (reset) begin
      data_901 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_901 <= data_900;
        end
      end
    end
    if (reset) begin
      data_902 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_902 <= data_901;
        end
      end
    end
    if (reset) begin
      data_903 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_903 <= data_902;
        end
      end
    end
    if (reset) begin
      data_904 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_904 <= data_903;
        end
      end
    end
    if (reset) begin
      data_905 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_905 <= data_904;
        end
      end
    end
    if (reset) begin
      data_906 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_906 <= data_905;
        end
      end
    end
    if (reset) begin
      data_907 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_907 <= data_906;
        end
      end
    end
    if (reset) begin
      data_908 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_908 <= data_907;
        end
      end
    end
    if (reset) begin
      data_909 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_909 <= data_908;
        end
      end
    end
    if (reset) begin
      data_910 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_910 <= data_909;
        end
      end
    end
    if (reset) begin
      data_911 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_911 <= data_910;
        end
      end
    end
    if (reset) begin
      data_912 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_912 <= data_911;
        end
      end
    end
    if (reset) begin
      data_913 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_913 <= data_912;
        end
      end
    end
    if (reset) begin
      data_914 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_914 <= data_913;
        end
      end
    end
    if (reset) begin
      data_915 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_915 <= data_914;
        end
      end
    end
    if (reset) begin
      data_916 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_916 <= data_915;
        end
      end
    end
    if (reset) begin
      data_917 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_917 <= data_916;
        end
      end
    end
    if (reset) begin
      data_918 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_918 <= data_917;
        end
      end
    end
    if (reset) begin
      data_919 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_919 <= data_918;
        end
      end
    end
    if (reset) begin
      data_920 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_920 <= data_919;
        end
      end
    end
    if (reset) begin
      data_921 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_921 <= data_920;
        end
      end
    end
    if (reset) begin
      data_922 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_922 <= data_921;
        end
      end
    end
    if (reset) begin
      data_923 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_923 <= data_922;
        end
      end
    end
    if (reset) begin
      data_924 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_924 <= data_923;
        end
      end
    end
    if (reset) begin
      data_925 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_925 <= data_924;
        end
      end
    end
    if (reset) begin
      data_926 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_926 <= data_925;
        end
      end
    end
    if (reset) begin
      data_927 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_927 <= data_926;
        end
      end
    end
    if (reset) begin
      data_928 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_928 <= data_927;
        end
      end
    end
    if (reset) begin
      data_929 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_929 <= data_928;
        end
      end
    end
    if (reset) begin
      data_930 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_930 <= data_929;
        end
      end
    end
    if (reset) begin
      data_931 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_931 <= data_930;
        end
      end
    end
    if (reset) begin
      data_932 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_932 <= data_931;
        end
      end
    end
    if (reset) begin
      data_933 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_933 <= data_932;
        end
      end
    end
    if (reset) begin
      data_934 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_934 <= data_933;
        end
      end
    end
    if (reset) begin
      data_935 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_935 <= data_934;
        end
      end
    end
    if (reset) begin
      data_936 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_936 <= data_935;
        end
      end
    end
    if (reset) begin
      data_937 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_937 <= data_936;
        end
      end
    end
    if (reset) begin
      data_938 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_938 <= data_937;
        end
      end
    end
    if (reset) begin
      data_939 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_939 <= data_938;
        end
      end
    end
    if (reset) begin
      data_940 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_940 <= data_939;
        end
      end
    end
    if (reset) begin
      data_941 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_941 <= data_940;
        end
      end
    end
    if (reset) begin
      data_942 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_942 <= data_941;
        end
      end
    end
    if (reset) begin
      data_943 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_943 <= data_942;
        end
      end
    end
    if (reset) begin
      data_944 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_944 <= data_943;
        end
      end
    end
    if (reset) begin
      data_945 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_945 <= data_944;
        end
      end
    end
    if (reset) begin
      data_946 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_946 <= data_945;
        end
      end
    end
    if (reset) begin
      data_947 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_947 <= data_946;
        end
      end
    end
    if (reset) begin
      data_948 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_948 <= data_947;
        end
      end
    end
    if (reset) begin
      data_949 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_949 <= data_948;
        end
      end
    end
    if (reset) begin
      data_950 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_950 <= data_949;
        end
      end
    end
    if (reset) begin
      data_951 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_951 <= data_950;
        end
      end
    end
    if (reset) begin
      data_952 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_952 <= data_951;
        end
      end
    end
    if (reset) begin
      data_953 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_953 <= data_952;
        end
      end
    end
    if (reset) begin
      data_954 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_954 <= data_953;
        end
      end
    end
    if (reset) begin
      data_955 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_955 <= data_954;
        end
      end
    end
    if (reset) begin
      data_956 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_956 <= data_955;
        end
      end
    end
    if (reset) begin
      data_957 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_957 <= data_956;
        end
      end
    end
    if (reset) begin
      data_958 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_958 <= data_957;
        end
      end
    end
    if (reset) begin
      data_959 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_959 <= data_958;
        end
      end
    end
    if (reset) begin
      data_960 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_960 <= data_959;
        end
      end
    end
    if (reset) begin
      data_961 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_961 <= data_960;
        end
      end
    end
    if (reset) begin
      data_962 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_962 <= data_961;
        end
      end
    end
    if (reset) begin
      data_963 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_963 <= data_962;
        end
      end
    end
    if (reset) begin
      data_964 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_964 <= data_963;
        end
      end
    end
    if (reset) begin
      data_965 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_965 <= data_964;
        end
      end
    end
    if (reset) begin
      data_966 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_966 <= data_965;
        end
      end
    end
    if (reset) begin
      data_967 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_967 <= data_966;
        end
      end
    end
    if (reset) begin
      data_968 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_968 <= data_967;
        end
      end
    end
    if (reset) begin
      data_969 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_969 <= data_968;
        end
      end
    end
    if (reset) begin
      data_970 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_970 <= data_969;
        end
      end
    end
    if (reset) begin
      data_971 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_971 <= data_970;
        end
      end
    end
    if (reset) begin
      data_972 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_972 <= data_971;
        end
      end
    end
    if (reset) begin
      data_973 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_973 <= data_972;
        end
      end
    end
    if (reset) begin
      data_974 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_974 <= data_973;
        end
      end
    end
    if (reset) begin
      data_975 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_975 <= data_974;
        end
      end
    end
    if (reset) begin
      data_976 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_976 <= data_975;
        end
      end
    end
    if (reset) begin
      data_977 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_977 <= data_976;
        end
      end
    end
    if (reset) begin
      data_978 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_978 <= data_977;
        end
      end
    end
    if (reset) begin
      data_979 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_979 <= data_978;
        end
      end
    end
    if (reset) begin
      data_980 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_980 <= data_979;
        end
      end
    end
    if (reset) begin
      data_981 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_981 <= data_980;
        end
      end
    end
    if (reset) begin
      data_982 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_982 <= data_981;
        end
      end
    end
    if (reset) begin
      data_983 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_983 <= data_982;
        end
      end
    end
    if (reset) begin
      data_984 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_984 <= data_983;
        end
      end
    end
    if (reset) begin
      data_985 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_985 <= data_984;
        end
      end
    end
    if (reset) begin
      data_986 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_986 <= data_985;
        end
      end
    end
    if (reset) begin
      data_987 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_987 <= data_986;
        end
      end
    end
    if (reset) begin
      data_988 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_988 <= data_987;
        end
      end
    end
    if (reset) begin
      data_989 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_989 <= data_988;
        end
      end
    end
    if (reset) begin
      data_990 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_990 <= data_989;
        end
      end
    end
    if (reset) begin
      data_991 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_991 <= data_990;
        end
      end
    end
    if (reset) begin
      data_992 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_992 <= data_991;
        end
      end
    end
    if (reset) begin
      data_993 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_993 <= data_992;
        end
      end
    end
    if (reset) begin
      data_994 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_994 <= data_993;
        end
      end
    end
    if (reset) begin
      data_995 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_995 <= data_994;
        end
      end
    end
    if (reset) begin
      data_996 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_996 <= data_995;
        end
      end
    end
    if (reset) begin
      data_997 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_997 <= data_996;
        end
      end
    end
    if (reset) begin
      data_998 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_998 <= data_997;
        end
      end
    end
    if (reset) begin
      data_999 <= 32'h0;
    end else if (valid) begin
      if (!(insn[6:0] == 7'hb)) begin
        if (insn[6:0] == 7'h2b) begin
          data_999 <= data_998;
        end
      end
    end
    if (reset) begin
      result <= 64'h0;
    end else if (valid) begin
      if (insn[6:0] == 7'hb) begin
        result <= {{32'd0}, _GEN_1999};
      end else if (insn[6:0] == 7'h2b) begin
        result <= {{32'd0}, data_0};
      end else begin
        result <= _GEN_2000;
      end
    end
  end
endmodule
