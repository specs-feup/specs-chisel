module TestDataMirror(
  input   clock,
  input   reset
);
endmodule
